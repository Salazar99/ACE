`timescale 1ns/1ns

module test;

  // Import the simplified package for ALU operations and parameters.
  import ibex_pkg::*;

  // Testbench parameters
  localparam CLK_PERIOD = 10; // 10 ns clock period

  // DUT signals
  logic clk;
  logic rst_n;
  alu_op_e operator_i;
  logic [31:0] operand_a_i;
  logic [31:0] operand_b_i;
  logic instr_first_cycle_i;
  logic [32:0] multdiv_operand_a_i;
  logic [32:0] multdiv_operand_b_i;
  logic multdiv_sel_i;
  logic [31:0] imd_val_q_i [2];
  logic [31:0] imd_val_d_o [2];
  logic [1:0] imd_val_we_o;
  logic [31:0] adder_result_o;
  logic [33:0] adder_result_ext_o;
  logic [31:0] result_o;
  logic comparison_result_o;
  logic is_equal_result_o;

  // Instantiate the Device Under Test (DUT)
  ibex_alu #(.RV32B(RV32BFull))
  i_ibex_alu (
    .operator_i          (operator_i),
    .operand_a_i         (operand_a_i),
    .operand_b_i         (operand_b_i),
    .instr_first_cycle_i (instr_first_cycle_i),
    .multdiv_operand_a_i (multdiv_operand_a_i),
    .multdiv_operand_b_i (multdiv_operand_b_i),
    .multdiv_sel_i       (multdiv_sel_i),
    .imd_val_q_i         (imd_val_q_i),
    .imd_val_d_o         (imd_val_d_o),
    .imd_val_we_o        (imd_val_we_o),
    .adder_result_o      (adder_result_o),
    .adder_result_ext_o  (adder_result_ext_o),
    .result_o            (result_o),
    .comparison_result_o (comparison_result_o),
    .is_equal_result_o   (is_equal_result_o)
  );


  always #5 clk = ~clk;


  initial begin

    $dumpfile("ibex_alu_1.vcd");

    $dumpvars(0, test);

    clk = 0;

    rst_n = 1;

    operator_i = ALU_SUB;

    operand_a_i = 7;

    operand_b_i = 1;

    #10;

    operand_a_i = 2;

    operand_b_i = 13;

    #10;

    operand_a_i = 17;

    operand_b_i = 20;

    #10;

    operand_a_i = 7;

    operand_b_i = 12;

    #10;

    operand_a_i = 11;

    operand_b_i = 9;

    #10;

    operand_a_i = 19;

    operand_b_i = 20;

    #10;

    operand_a_i = 16;

    operand_b_i = 4;

    #10;

    operand_a_i = 1;

    operand_b_i = 10;

    #10;

    operand_a_i = 9;

    operand_b_i = 15;

    #10;

    operand_a_i = 20;

    operand_b_i = 11;

    #10;

    operand_a_i = 19;

    operand_b_i = 13;

    #10;

    operand_a_i = 8;

    operand_b_i = 9;

    #10;

    operand_a_i = 11;

    operand_b_i = 7;

    #10;

    operand_a_i = 3;

    operand_b_i = 12;

    #10;

    operand_a_i = 2;

    operand_b_i = 12;

    #10;

    operand_a_i = 19;

    operand_b_i = 16;

    #10;

    operand_a_i = 15;

    operand_b_i = 9;

    #10;

    operand_a_i = 3;

    operand_b_i = 20;

    #10;

    operand_a_i = 19;

    operand_b_i = 4;

    #10;

    operand_a_i = 9;

    operand_b_i = 13;

    #10;

    operand_a_i = 7;

    operand_b_i = 20;

    #10;

    operand_a_i = 4;

    operand_b_i = 19;

    #10;

    operand_a_i = 10;

    operand_b_i = 16;

    #10;

    operand_a_i = 13;

    operand_b_i = 6;

    #10;

    operand_a_i = 20;

    operand_b_i = 8;

    #10;

    operand_a_i = 6;

    operand_b_i = 4;

    #10;

    operand_a_i = 10;

    operand_b_i = 6;

    #10;

    operand_a_i = 15;

    operand_b_i = 11;

    #10;

    operand_a_i = 5;

    operand_b_i = 6;

    #10;

    operand_a_i = 17;

    operand_b_i = 9;

    #10;

    operand_a_i = 14;

    operand_b_i = 19;

    #10;

    operand_a_i = 5;

    operand_b_i = 19;

    #10;

    operand_a_i = 18;

    operand_b_i = 9;

    #10;

    operand_a_i = 6;

    operand_b_i = 15;

    #10;

    operand_a_i = 1;

    operand_b_i = 3;

    #10;

    operand_a_i = 8;

    operand_b_i = 4;

    #10;

    operand_a_i = 9;

    operand_b_i = 19;

    #10;

    operand_a_i = 19;

    operand_b_i = 8;

    #10;

    operand_a_i = 10;

    operand_b_i = 8;

    #10;

    operand_a_i = 10;

    operand_b_i = 17;

    #10;

    operand_a_i = 10;

    operand_b_i = 11;

    #10;

    operand_a_i = 3;

    operand_b_i = 4;

    #10;

    operand_a_i = 12;

    operand_b_i = 1;

    #10;

    operand_a_i = 19;

    operand_b_i = 2;

    #10;

    operand_a_i = 3;

    operand_b_i = 16;

    #10;

    operand_a_i = 3;

    operand_b_i = 5;

    #10;

    operand_a_i = 11;

    operand_b_i = 15;

    #10;

    operand_a_i = 11;

    operand_b_i = 10;

    #10;

    operand_a_i = 1;

    operand_b_i = 6;

    #10;

    operand_a_i = 18;

    operand_b_i = 2;

    #10;

    operand_a_i = 12;

    operand_b_i = 3;

    #10;

    operand_a_i = 2;

    operand_b_i = 16;

    #10;

    operand_a_i = 4;

    operand_b_i = 16;

    #10;

    operand_a_i = 9;

    operand_b_i = 19;

    #10;

    operand_a_i = 14;

    operand_b_i = 9;

    #10;

    operand_a_i = 12;

    operand_b_i = 3;

    #10;

    operand_a_i = 17;

    operand_b_i = 4;

    #10;

    operand_a_i = 17;

    operand_b_i = 15;

    #10;

    operand_a_i = 8;

    operand_b_i = 18;

    #10;

    operand_a_i = 15;

    operand_b_i = 16;

    #10;

    operand_a_i = 14;

    operand_b_i = 4;

    #10;

    operand_a_i = 16;

    operand_b_i = 2;

    #10;

    operand_a_i = 20;

    operand_b_i = 1;

    #10;

    operand_a_i = 17;

    operand_b_i = 5;

    #10;

    operand_a_i = 17;

    operand_b_i = 16;

    #10;

    operand_a_i = 6;

    operand_b_i = 17;

    #10;

    operand_a_i = 4;

    operand_b_i = 13;

    #10;

    operand_a_i = 14;

    operand_b_i = 4;

    #10;

    operand_a_i = 16;

    operand_b_i = 1;

    #10;

    operand_a_i = 9;

    operand_b_i = 19;

    #10;

    operand_a_i = 6;

    operand_b_i = 8;

    #10;

    operand_a_i = 17;

    operand_b_i = 15;

    #10;

    operand_a_i = 11;

    operand_b_i = 2;

    #10;

    operand_a_i = 10;

    operand_b_i = 11;

    #10;

    operand_a_i = 17;

    operand_b_i = 14;

    #10;

    operand_a_i = 10;

    operand_b_i = 6;

    #10;

    operand_a_i = 6;

    operand_b_i = 15;

    #10;

    operand_a_i = 8;

    operand_b_i = 16;

    #10;

    operand_a_i = 6;

    operand_b_i = 13;

    #10;

    operand_a_i = 13;

    operand_b_i = 1;

    #10;

    operand_a_i = 18;

    operand_b_i = 9;

    #10;

    operand_a_i = 1;

    operand_b_i = 5;

    #10;

    operand_a_i = 5;

    operand_b_i = 4;

    #10;

    operand_a_i = 19;

    operand_b_i = 2;

    #10;

    operand_a_i = 20;

    operand_b_i = 16;

    #10;

    operand_a_i = 6;

    operand_b_i = 8;

    #10;

    operand_a_i = 10;

    operand_b_i = 15;

    #10;

    operand_a_i = 2;

    operand_b_i = 10;

    #10;

    operand_a_i = 9;

    operand_b_i = 7;

    #10;

    operand_a_i = 10;

    operand_b_i = 20;

    #10;

    operand_a_i = 2;

    operand_b_i = 17;

    #10;

    operand_a_i = 1;

    operand_b_i = 16;

    #10;

    operand_a_i = 11;

    operand_b_i = 3;

    #10;

    operand_a_i = 15;

    operand_b_i = 5;

    #10;

    operand_a_i = 8;

    operand_b_i = 15;

    #10;

    operand_a_i = 2;

    operand_b_i = 8;

    #10;

    operand_a_i = 18;

    operand_b_i = 1;

    #10;

    operand_a_i = 13;

    operand_b_i = 9;

    #10;

    operand_a_i = 13;

    operand_b_i = 1;

    #10;

    operand_a_i = 12;

    operand_b_i = 17;

    #10;

    operand_a_i = 14;

    operand_b_i = 6;

    #10;

    operand_a_i = 12;

    operand_b_i = 19;

    #10;

    operand_a_i = 5;

    operand_b_i = 7;

    #10;

    operand_a_i = 3;

    operand_b_i = 5;

    #10;

    operand_a_i = 7;

    operand_b_i = 6;

    #10;

    operand_a_i = 9;

    operand_b_i = 19;

    #10;

    operand_a_i = 1;

    operand_b_i = 7;

    #10;

    operand_a_i = 16;

    operand_b_i = 17;

    #10;

    operand_a_i = 16;

    operand_b_i = 8;

    #10;

    operand_a_i = 19;

    operand_b_i = 16;

    #10;

    operand_a_i = 6;

    operand_b_i = 16;

    #10;

    operand_a_i = 1;

    operand_b_i = 13;

    #10;

    operand_a_i = 19;

    operand_b_i = 16;

    #10;

    operand_a_i = 18;

    operand_b_i = 4;

    #10;

    operand_a_i = 1;

    operand_b_i = 5;

    #10;

    operand_a_i = 9;

    operand_b_i = 8;

    #10;

    operand_a_i = 11;

    operand_b_i = 14;

    #10;

    operand_a_i = 14;

    operand_b_i = 15;

    #10;

    operand_a_i = 15;

    operand_b_i = 17;

    #10;

    operand_a_i = 1;

    operand_b_i = 12;

    #10;

    operand_a_i = 10;

    operand_b_i = 6;

    #10;

    operand_a_i = 9;

    operand_b_i = 18;

    #10;

    operand_a_i = 5;

    operand_b_i = 19;

    #10;

    operand_a_i = 8;

    operand_b_i = 11;

    #10;

    operand_a_i = 7;

    operand_b_i = 18;

    #10;

    operand_a_i = 8;

    operand_b_i = 16;

    #10;

    operand_a_i = 13;

    operand_b_i = 8;

    #10;

    operand_a_i = 1;

    operand_b_i = 16;

    #10;

    operand_a_i = 7;

    operand_b_i = 20;

    #10;

    operand_a_i = 1;

    operand_b_i = 11;

    #10;

    operand_a_i = 15;

    operand_b_i = 9;

    #10;

    operand_a_i = 13;

    operand_b_i = 17;

    #10;

    operand_a_i = 14;

    operand_b_i = 16;

    #10;

    operand_a_i = 17;

    operand_b_i = 15;

    #10;

    operand_a_i = 2;

    operand_b_i = 10;

    #10;

    operand_a_i = 14;

    operand_b_i = 13;

    #10;

    operand_a_i = 11;

    operand_b_i = 10;

    #10;

    operand_a_i = 2;

    operand_b_i = 8;

    #10;

    operand_a_i = 11;

    operand_b_i = 4;

    #10;

    operand_a_i = 18;

    operand_b_i = 13;

    #10;

    operand_a_i = 4;

    operand_b_i = 7;

    #10;

    operand_a_i = 16;

    operand_b_i = 3;

    #10;

    operand_a_i = 7;

    operand_b_i = 18;

    #10;

    operand_a_i = 12;

    operand_b_i = 4;

    #10;

    operand_a_i = 6;

    operand_b_i = 4;

    #10;

    operand_a_i = 9;

    operand_b_i = 6;

    #10;

    operand_a_i = 14;

    operand_b_i = 1;

    #10;

    operand_a_i = 1;

    operand_b_i = 15;

    #10;

    operand_a_i = 20;

    operand_b_i = 8;

    #10;

    operand_a_i = 20;

    operand_b_i = 1;

    #10;

    operand_a_i = 17;

    operand_b_i = 4;

    #10;

    operand_a_i = 12;

    operand_b_i = 4;

    #10;

    operand_a_i = 17;

    operand_b_i = 9;

    #10;

    operand_a_i = 11;

    operand_b_i = 7;

    #10;

    operand_a_i = 4;

    operand_b_i = 16;

    #10;

    operand_a_i = 10;

    operand_b_i = 9;

    #10;

    operand_a_i = 8;

    operand_b_i = 18;

    #10;

    operand_a_i = 10;

    operand_b_i = 11;

    #10;

    operand_a_i = 6;

    operand_b_i = 1;

    #10;

    operand_a_i = 3;

    operand_b_i = 14;

    #10;

    operand_a_i = 10;

    operand_b_i = 9;

    #10;

    operand_a_i = 16;

    operand_b_i = 2;

    #10;

    operand_a_i = 4;

    operand_b_i = 9;

    #10;

    operand_a_i = 10;

    operand_b_i = 19;

    #10;

    operand_a_i = 3;

    operand_b_i = 20;

    #10;

    operand_a_i = 2;

    operand_b_i = 10;

    #10;

    operand_a_i = 13;

    operand_b_i = 6;

    #10;

    operand_a_i = 14;

    operand_b_i = 5;

    #10;

    operand_a_i = 19;

    operand_b_i = 2;

    #10;

    operand_a_i = 13;

    operand_b_i = 14;

    #10;

    operand_a_i = 2;

    operand_b_i = 7;

    #10;

    operand_a_i = 13;

    operand_b_i = 2;

    #10;

    operand_a_i = 6;

    operand_b_i = 16;

    #10;

    operand_a_i = 6;

    operand_b_i = 14;

    #10;

    operand_a_i = 5;

    operand_b_i = 7;

    #10;

    operand_a_i = 15;

    operand_b_i = 4;

    #10;

    operand_a_i = 11;

    operand_b_i = 19;

    #10;

    operand_a_i = 12;

    operand_b_i = 11;

    #10;

    operand_a_i = 7;

    operand_b_i = 10;

    #10;

    operand_a_i = 14;

    operand_b_i = 17;

    #10;

    operand_a_i = 19;

    operand_b_i = 5;

    #10;

    operand_a_i = 2;

    operand_b_i = 14;

    #10;

    operand_a_i = 9;

    operand_b_i = 20;

    #10;

    operand_a_i = 13;

    operand_b_i = 5;

    #10;

    operand_a_i = 8;

    operand_b_i = 18;

    #10;

    operand_a_i = 9;

    operand_b_i = 20;

    #10;

    operand_a_i = 1;

    operand_b_i = 11;

    #10;

    operand_a_i = 17;

    operand_b_i = 16;

    #10;

    operand_a_i = 14;

    operand_b_i = 11;

    #10;

    operand_a_i = 4;

    operand_b_i = 13;

    #10;

    operand_a_i = 5;

    operand_b_i = 17;

    #10;

    operand_a_i = 17;

    operand_b_i = 15;

    #10;

    operand_a_i = 12;

    operand_b_i = 5;

    #10;

    operand_a_i = 18;

    operand_b_i = 3;

    #10;

    operand_a_i = 6;

    operand_b_i = 16;

    #10;

    operand_a_i = 15;

    operand_b_i = 20;

    #10;

    operand_a_i = 18;

    operand_b_i = 3;

    #10;

    operand_a_i = 2;

    operand_b_i = 6;

    #10;

    operand_a_i = 14;

    operand_b_i = 4;

    #10;

    operand_a_i = 11;

    operand_b_i = 20;

    #10;

    operand_a_i = 7;

    operand_b_i = 3;

    #10;

    operand_a_i = 20;

    operand_b_i = 13;

    #10;

    operand_a_i = 18;

    operand_b_i = 19;

    #10;

    operand_a_i = 9;

    operand_b_i = 8;

    #10;

    operand_a_i = 11;

    operand_b_i = 3;

    #10;

    operand_a_i = 14;

    operand_b_i = 15;

    #10;

    operand_a_i = 7;

    operand_b_i = 9;

    #10;

    operand_a_i = 14;

    operand_b_i = 17;

    #10;

    operand_a_i = 3;

    operand_b_i = 15;

    #10;

    operand_a_i = 6;

    operand_b_i = 19;

    #10;

    operand_a_i = 20;

    operand_b_i = 5;

    #10;

    operand_a_i = 17;

    operand_b_i = 19;

    #10;

    operand_a_i = 6;

    operand_b_i = 13;

    #10;

    operand_a_i = 8;

    operand_b_i = 4;

    #10;

    operand_a_i = 11;

    operand_b_i = 13;

    #10;

    operand_a_i = 16;

    operand_b_i = 18;

    #10;

    operand_a_i = 10;

    operand_b_i = 19;

    #10;

    operand_a_i = 11;

    operand_b_i = 20;

    #10;

    operand_a_i = 10;

    operand_b_i = 15;

    #10;

    operand_a_i = 14;

    operand_b_i = 17;

    #10;

    operand_a_i = 7;

    operand_b_i = 17;

    #10;

    operand_a_i = 9;

    operand_b_i = 17;

    #10;

    operand_a_i = 7;

    operand_b_i = 8;

    #10;

    operand_a_i = 9;

    operand_b_i = 2;

    #10;

    operand_a_i = 19;

    operand_b_i = 18;

    #10;

    operand_a_i = 5;

    operand_b_i = 17;

    #10;

    operand_a_i = 2;

    operand_b_i = 14;

    #10;

    operand_a_i = 20;

    operand_b_i = 12;

    #10;

    operand_a_i = 2;

    operand_b_i = 12;

    #10;

    operand_a_i = 17;

    operand_b_i = 3;

    #10;

    operand_a_i = 4;

    operand_b_i = 13;

    #10;

    operand_a_i = 12;

    operand_b_i = 20;

    #10;

    operand_a_i = 18;

    operand_b_i = 12;

    #10;

    operand_a_i = 6;

    operand_b_i = 7;

    #10;

    operand_a_i = 7;

    operand_b_i = 2;

    #10;

    operand_a_i = 5;

    operand_b_i = 9;

    #10;

    operand_a_i = 14;

    operand_b_i = 18;

    #10;

    operand_a_i = 6;

    operand_b_i = 5;

    #10;

    operand_a_i = 11;

    operand_b_i = 9;

    #10;

    operand_a_i = 13;

    operand_b_i = 4;

    #10;

    operand_a_i = 17;

    operand_b_i = 1;

    #10;

    operand_a_i = 6;

    operand_b_i = 1;

    #10;

    operand_a_i = 19;

    operand_b_i = 9;

    #10;

    operand_a_i = 9;

    operand_b_i = 17;

    #10;

    operand_a_i = 18;

    operand_b_i = 10;

    #10;

    operand_a_i = 16;

    operand_b_i = 9;

    #10;

    operand_a_i = 14;

    operand_b_i = 13;

    #10;

    operand_a_i = 16;

    operand_b_i = 6;

    #10;

    operand_a_i = 14;

    operand_b_i = 20;

    #10;

    operand_a_i = 17;

    operand_b_i = 19;

    #10;

    operand_a_i = 7;

    operand_b_i = 6;

    #10;

    operand_a_i = 10;

    operand_b_i = 12;

    #10;

    operand_a_i = 12;

    operand_b_i = 15;

    #10;

    operand_a_i = 15;

    operand_b_i = 7;

    #10;

    operand_a_i = 17;

    operand_b_i = 13;

    #10;

    operand_a_i = 10;

    operand_b_i = 14;

    #10;

    operand_a_i = 20;

    operand_b_i = 18;

    #10;

    operand_a_i = 17;

    operand_b_i = 8;

    #10;

    operand_a_i = 4;

    operand_b_i = 3;

    #10;

    operand_a_i = 7;

    operand_b_i = 14;

    #10;

    operand_a_i = 10;

    operand_b_i = 19;

    #10;

    operand_a_i = 13;

    operand_b_i = 14;

    #10;

    operand_a_i = 20;

    operand_b_i = 2;

    #10;

    operand_a_i = 10;

    operand_b_i = 5;

    #10;

    operand_a_i = 9;

    operand_b_i = 10;

    #10;

    operand_a_i = 2;

    operand_b_i = 19;

    #10;

    operand_a_i = 18;

    operand_b_i = 10;

    #10;

    operand_a_i = 12;

    operand_b_i = 14;

    #10;

    operand_a_i = 20;

    operand_b_i = 11;

    #10;

    operand_a_i = 4;

    operand_b_i = 3;

    #10;

    operand_a_i = 1;

    operand_b_i = 15;

    #10;

    operand_a_i = 3;

    operand_b_i = 7;

    #10;

    operand_a_i = 5;

    operand_b_i = 20;

    #10;

    operand_a_i = 9;

    operand_b_i = 15;

    #10;

    operand_a_i = 17;

    operand_b_i = 10;

    #10;

    operand_a_i = 14;

    operand_b_i = 18;

    #10;

    operand_a_i = 2;

    operand_b_i = 9;

    #10;

    operand_a_i = 3;

    operand_b_i = 6;

    #10;

    operand_a_i = 3;

    operand_b_i = 11;

    #10;

    operand_a_i = 8;

    operand_b_i = 20;

    #10;

    operand_a_i = 16;

    operand_b_i = 15;

    #10;

    operand_a_i = 9;

    operand_b_i = 7;

    #10;

    operand_a_i = 12;

    operand_b_i = 15;

    #10;

    operand_a_i = 17;

    operand_b_i = 9;

    #10;

    operand_a_i = 6;

    operand_b_i = 14;

    #10;

    operand_a_i = 11;

    operand_b_i = 19;

    #10;

    operand_a_i = 8;

    operand_b_i = 2;

    #10;

    operand_a_i = 15;

    operand_b_i = 10;

    #10;

    operand_a_i = 3;

    operand_b_i = 17;

    #10;

    operand_a_i = 13;

    operand_b_i = 19;

    #10;

    operand_a_i = 11;

    operand_b_i = 13;

    #10;

    operand_a_i = 8;

    operand_b_i = 16;

    #10;

    operand_a_i = 15;

    operand_b_i = 1;

    #10;

    operand_a_i = 7;

    operand_b_i = 6;

    #10;

    operand_a_i = 7;

    operand_b_i = 18;

    #10;

    operand_a_i = 8;

    operand_b_i = 16;

    #10;

    operand_a_i = 16;

    operand_b_i = 7;

    #10;

    operand_a_i = 2;

    operand_b_i = 14;

    #10;

    operand_a_i = 1;

    operand_b_i = 17;

    #10;

    operand_a_i = 8;

    operand_b_i = 2;

    #10;

    operand_a_i = 16;

    operand_b_i = 11;

    #10;

    operand_a_i = 20;

    operand_b_i = 4;

    #10;

    operand_a_i = 10;

    operand_b_i = 3;

    #10;

    operand_a_i = 19;

    operand_b_i = 4;

    #10;

    operand_a_i = 1;

    operand_b_i = 12;

    #10;

    operand_a_i = 12;

    operand_b_i = 19;

    #10;

    operand_a_i = 1;

    operand_b_i = 10;

    #10;

    operand_a_i = 7;

    operand_b_i = 14;

    #10;

    operand_a_i = 20;

    operand_b_i = 9;

    #10;

    operand_a_i = 20;

    operand_b_i = 4;

    #10;

    operand_a_i = 8;

    operand_b_i = 13;

    #10;

    operand_a_i = 12;

    operand_b_i = 11;

    #10;

    operand_a_i = 9;

    operand_b_i = 10;

    #10;

    operand_a_i = 6;

    operand_b_i = 7;

    #10;

    operand_a_i = 2;

    operand_b_i = 15;

    #10;

    operand_a_i = 20;

    operand_b_i = 1;

    #10;

    operand_a_i = 4;

    operand_b_i = 20;

    #10;

    operand_a_i = 15;

    operand_b_i = 14;

    #10;

    operand_a_i = 14;

    operand_b_i = 18;

    #10;

    operand_a_i = 1;

    operand_b_i = 20;

    #10;

    operand_a_i = 11;

    operand_b_i = 12;

    #10;

    operand_a_i = 5;

    operand_b_i = 6;

    #10;

    operand_a_i = 13;

    operand_b_i = 14;

    #10;

    operand_a_i = 1;

    operand_b_i = 10;

    #10;

    operand_a_i = 7;

    operand_b_i = 11;

    #10;

    operand_a_i = 7;

    operand_b_i = 15;

    #10;

    operand_a_i = 3;

    operand_b_i = 14;

    #10;

    operand_a_i = 16;

    operand_b_i = 13;

    #10;

    operand_a_i = 14;

    operand_b_i = 5;

    #10;

    operand_a_i = 18;

    operand_b_i = 16;

    #10;

    operand_a_i = 19;

    operand_b_i = 14;

    #10;

    operand_a_i = 6;

    operand_b_i = 11;

    #10;

    operand_a_i = 11;

    operand_b_i = 12;

    #10;

    operand_a_i = 6;

    operand_b_i = 8;

    #10;

    operand_a_i = 1;

    operand_b_i = 9;

    #10;

    operand_a_i = 7;

    operand_b_i = 18;

    #10;

    operand_a_i = 13;

    operand_b_i = 4;

    #10;

    operand_a_i = 4;

    operand_b_i = 8;

    #10;

    operand_a_i = 11;

    operand_b_i = 2;

    #10;

    operand_a_i = 14;

    operand_b_i = 3;

    #10;

    operand_a_i = 7;

    operand_b_i = 20;

    #10;

    operand_a_i = 12;

    operand_b_i = 8;

    #10;

    operand_a_i = 8;

    operand_b_i = 16;

    #10;

    operand_a_i = 20;

    operand_b_i = 10;

    #10;

    operand_a_i = 11;

    operand_b_i = 5;

    #10;

    operand_a_i = 5;

    operand_b_i = 6;

    #10;

    operand_a_i = 7;

    operand_b_i = 6;

    #10;

    operand_a_i = 5;

    operand_b_i = 19;

    #10;

    operand_a_i = 19;

    operand_b_i = 14;

    #10;

    operand_a_i = 11;

    operand_b_i = 14;

    #10;

    operand_a_i = 2;

    operand_b_i = 11;

    #10;

    operand_a_i = 18;

    operand_b_i = 1;

    #10;

    operand_a_i = 19;

    operand_b_i = 9;

    #10;

    operand_a_i = 8;

    operand_b_i = 9;

    #10;

    operand_a_i = 10;

    operand_b_i = 20;

    #10;

    operand_a_i = 2;

    operand_b_i = 1;

    #10;

    operand_a_i = 4;

    operand_b_i = 6;

    #10;

    operand_a_i = 16;

    operand_b_i = 8;

    #10;

    operand_a_i = 6;

    operand_b_i = 19;

    #10;

    operand_a_i = 9;

    operand_b_i = 17;

    #10;

    operand_a_i = 19;

    operand_b_i = 11;

    #10;

    operand_a_i = 2;

    operand_b_i = 7;

    #10;

    operand_a_i = 6;

    operand_b_i = 8;

    #10;

    operand_a_i = 9;

    operand_b_i = 10;

    #10;

    operand_a_i = 8;

    operand_b_i = 15;

    #10;

    operand_a_i = 19;

    operand_b_i = 10;

    #10;

    operand_a_i = 15;

    operand_b_i = 16;

    #10;

    operand_a_i = 12;

    operand_b_i = 6;

    #10;

    operand_a_i = 19;

    operand_b_i = 12;

    #10;

    operand_a_i = 19;

    operand_b_i = 9;

    #10;

    operand_a_i = 13;

    operand_b_i = 10;

    #10;

    operand_a_i = 12;

    operand_b_i = 16;

    #10;

    operand_a_i = 5;

    operand_b_i = 14;

    #10;

    operand_a_i = 14;

    operand_b_i = 13;

    #10;

    operand_a_i = 2;

    operand_b_i = 16;

    #10;

    operand_a_i = 13;

    operand_b_i = 9;

    #10;

    operand_a_i = 2;

    operand_b_i = 3;

    #10;

    operand_a_i = 7;

    operand_b_i = 10;

    #10;

    operand_a_i = 3;

    operand_b_i = 16;

    #10;

    operand_a_i = 15;

    operand_b_i = 1;

    #10;

    operand_a_i = 18;

    operand_b_i = 2;

    #10;

    operand_a_i = 15;

    operand_b_i = 18;

    #10;

    operand_a_i = 5;

    operand_b_i = 3;

    #10;

    operand_a_i = 5;

    operand_b_i = 7;

    #10;

    operand_a_i = 8;

    operand_b_i = 4;

    #10;

    operand_a_i = 2;

    operand_b_i = 17;

    #10;

    operand_a_i = 1;

    operand_b_i = 6;

    #10;

    operand_a_i = 18;

    operand_b_i = 12;

    #10;

    operand_a_i = 7;

    operand_b_i = 3;

    #10;

    operand_a_i = 3;

    operand_b_i = 11;

    #10;

    operand_a_i = 12;

    operand_b_i = 19;

    #10;

    operand_a_i = 2;

    operand_b_i = 15;

    #10;

    operand_a_i = 19;

    operand_b_i = 17;

    #10;

    operand_a_i = 13;

    operand_b_i = 1;

    #10;

    operand_a_i = 14;

    operand_b_i = 1;

    #10;

    operand_a_i = 14;

    operand_b_i = 17;

    #10;

    operand_a_i = 11;

    operand_b_i = 20;

    #10;

    operand_a_i = 6;

    operand_b_i = 9;

    #10;

    operand_a_i = 14;

    operand_b_i = 16;

    #10;

    operand_a_i = 18;

    operand_b_i = 17;

    #10;

    operand_a_i = 9;

    operand_b_i = 7;

    #10;

    operand_a_i = 1;

    operand_b_i = 16;

    #10;

    operand_a_i = 15;

    operand_b_i = 8;

    #10;

    operand_a_i = 6;

    operand_b_i = 3;

    #10;

    operand_a_i = 14;

    operand_b_i = 8;

    #10;

    operand_a_i = 4;

    operand_b_i = 3;

    #10;

    operand_a_i = 7;

    operand_b_i = 20;

    #10;

    operand_a_i = 2;

    operand_b_i = 19;

    #10;

    operand_a_i = 13;

    operand_b_i = 3;

    #10;

    operand_a_i = 3;

    operand_b_i = 16;

    #10;

    operand_a_i = 19;

    operand_b_i = 13;

    #10;

    operand_a_i = 7;

    operand_b_i = 8;

    #10;

    operand_a_i = 14;

    operand_b_i = 7;

    #10;

    operand_a_i = 13;

    operand_b_i = 1;

    #10;

    operand_a_i = 19;

    operand_b_i = 3;

    #10;

    operand_a_i = 1;

    operand_b_i = 16;

    #10;

    operand_a_i = 11;

    operand_b_i = 16;

    #10;

    operand_a_i = 13;

    operand_b_i = 7;

    #10;

    operand_a_i = 12;

    operand_b_i = 10;

    #10;

    operand_a_i = 9;

    operand_b_i = 17;

    #10;

    operand_a_i = 4;

    operand_b_i = 8;

    #10;

    operand_a_i = 12;

    operand_b_i = 2;

    #10;

    operand_a_i = 16;

    operand_b_i = 17;

    #10;

    operand_a_i = 5;

    operand_b_i = 14;

    #10;

    operand_a_i = 12;

    operand_b_i = 11;

    #10;

    operand_a_i = 9;

    operand_b_i = 7;

    #10;

    operand_a_i = 11;

    operand_b_i = 20;

    #10;

    operand_a_i = 12;

    operand_b_i = 19;

    #10;

    operand_a_i = 9;

    operand_b_i = 2;

    #10;

    operand_a_i = 20;

    operand_b_i = 11;

    #10;

    operand_a_i = 9;

    operand_b_i = 11;

    #10;

    operand_a_i = 15;

    operand_b_i = 1;

    #10;

    operand_a_i = 13;

    operand_b_i = 16;

    #10;

    operand_a_i = 11;

    operand_b_i = 7;

    #10;

    operand_a_i = 10;

    operand_b_i = 5;

    #10;

    operand_a_i = 10;

    operand_b_i = 2;

    #10;

    operand_a_i = 16;

    operand_b_i = 18;

    #10;

    operand_a_i = 15;

    operand_b_i = 12;

    #10;

    operand_a_i = 16;

    operand_b_i = 10;

    #10;

    operand_a_i = 16;

    operand_b_i = 20;

    #10;

    operand_a_i = 14;

    operand_b_i = 10;

    #10;

    operand_a_i = 16;

    operand_b_i = 7;

    #10;

    operand_a_i = 20;

    operand_b_i = 13;

    #10;

    operand_a_i = 19;

    operand_b_i = 9;

    #10;

    operand_a_i = 20;

    operand_b_i = 13;

    #10;

    operand_a_i = 12;

    operand_b_i = 15;

    #10;

    operand_a_i = 2;

    operand_b_i = 16;

    #10;

    operand_a_i = 17;

    operand_b_i = 11;

    #10;

    operand_a_i = 14;

    operand_b_i = 13;

    #10;

    operand_a_i = 6;

    operand_b_i = 8;

    #10;

    operand_a_i = 8;

    operand_b_i = 19;

    #10;

    operand_a_i = 2;

    operand_b_i = 1;

    #10;

    operand_a_i = 16;

    operand_b_i = 8;

    #10;

    operand_a_i = 16;

    operand_b_i = 17;

    #10;

    operand_a_i = 1;

    operand_b_i = 10;

    #10;

    operand_a_i = 8;

    operand_b_i = 16;

    #10;

    operand_a_i = 9;

    operand_b_i = 4;

    #10;

    operand_a_i = 17;

    operand_b_i = 3;

    #10;

    operand_a_i = 11;

    operand_b_i = 6;

    #10;

    operand_a_i = 14;

    operand_b_i = 8;

    #10;

    operand_a_i = 11;

    operand_b_i = 5;

    #10;

    operand_a_i = 1;

    operand_b_i = 20;

    #10;

    operand_a_i = 18;

    operand_b_i = 2;

    #10;

    operand_a_i = 16;

    operand_b_i = 8;

    #10;

    operand_a_i = 10;

    operand_b_i = 8;

    #10;

    operand_a_i = 11;

    operand_b_i = 20;

    #10;

    operand_a_i = 4;

    operand_b_i = 17;

    #10;

    operand_a_i = 19;

    operand_b_i = 11;

    #10;

    operand_a_i = 4;

    operand_b_i = 5;

    #10;

    operand_a_i = 14;

    operand_b_i = 11;

    #10;

    operand_a_i = 17;

    operand_b_i = 16;

    #10;

    operand_a_i = 13;

    operand_b_i = 8;

    #10;

    operand_a_i = 20;

    operand_b_i = 10;

    #10;

    operand_a_i = 10;

    operand_b_i = 15;

    #10;

    operand_a_i = 7;

    operand_b_i = 1;

    #10;

    operand_a_i = 14;

    operand_b_i = 7;

    #10;

    operand_a_i = 12;

    operand_b_i = 17;

    #10;

    operand_a_i = 5;

    operand_b_i = 2;

    #10;

    operand_a_i = 20;

    operand_b_i = 6;

    #10;

    operand_a_i = 2;

    operand_b_i = 3;

    #10;

    operand_a_i = 18;

    operand_b_i = 1;

    #10;

    operand_a_i = 17;

    operand_b_i = 15;

    #10;

    operand_a_i = 6;

    operand_b_i = 12;

    #10;

    operand_a_i = 15;

    operand_b_i = 11;

    #10;

    operand_a_i = 7;

    operand_b_i = 4;

    #10;

    operand_a_i = 9;

    operand_b_i = 15;

    #10;

    operand_a_i = 17;

    operand_b_i = 11;

    #10;

    operand_a_i = 1;

    operand_b_i = 8;

    #10;

    operand_a_i = 3;

    operand_b_i = 16;

    #10;

    operand_a_i = 9;

    operand_b_i = 11;

    #10;

    operand_a_i = 14;

    operand_b_i = 16;

    #10;

    operand_a_i = 9;

    operand_b_i = 3;

    #10;

    operand_a_i = 8;

    operand_b_i = 18;

    #10;

    operand_a_i = 4;

    operand_b_i = 8;

    #10;

    operand_a_i = 6;

    operand_b_i = 8;

    #10;

    operand_a_i = 16;

    operand_b_i = 10;

    #10;

    operand_a_i = 14;

    operand_b_i = 5;

    #10;

    operand_a_i = 12;

    operand_b_i = 6;

    #10;

    operand_a_i = 2;

    operand_b_i = 18;

    #10;

    operand_a_i = 4;

    operand_b_i = 11;

    #10;

    operand_a_i = 8;

    operand_b_i = 10;

    #10;

    operand_a_i = 1;

    operand_b_i = 10;

    #10;

    operand_a_i = 14;

    operand_b_i = 2;

    #10;

    operand_a_i = 1;

    operand_b_i = 19;

    #10;

    operand_a_i = 6;

    operand_b_i = 13;

    #10;

    operand_a_i = 3;

    operand_b_i = 6;

    #10;

    operand_a_i = 17;

    operand_b_i = 20;

    #10;

    operand_a_i = 12;

    operand_b_i = 15;

    #10;

    operand_a_i = 19;

    operand_b_i = 4;

    #10;

    operand_a_i = 8;

    operand_b_i = 7;

    #10;

    operand_a_i = 2;

    operand_b_i = 15;

    #10;

    operand_a_i = 13;

    operand_b_i = 15;

    #10;

    operand_a_i = 16;

    operand_b_i = 17;

    #10;

    operand_a_i = 6;

    operand_b_i = 17;

    #10;

    operand_a_i = 15;

    operand_b_i = 8;

    #10;

    operand_a_i = 13;

    operand_b_i = 11;

    #10;

    operand_a_i = 9;

    operand_b_i = 1;

    #10;

    operand_a_i = 8;

    operand_b_i = 17;

    #10;

    operand_a_i = 9;

    operand_b_i = 20;

    #10;

    operand_a_i = 6;

    operand_b_i = 4;

    #10;

    operand_a_i = 6;

    operand_b_i = 1;

    #10;

    operand_a_i = 8;

    operand_b_i = 13;

    #10;

    operand_a_i = 6;

    operand_b_i = 12;

    #10;

    operand_a_i = 7;

    operand_b_i = 14;

    #10;

    operand_a_i = 19;

    operand_b_i = 16;

    #10;

    operand_a_i = 16;

    operand_b_i = 14;

    #10;

    operand_a_i = 20;

    operand_b_i = 5;

    #10;

    operand_a_i = 2;

    operand_b_i = 11;

    #10;

    operand_a_i = 2;

    operand_b_i = 8;

    #10;

    operand_a_i = 8;

    operand_b_i = 10;

    #10;

    operand_a_i = 19;

    operand_b_i = 15;

    #10;

    operand_a_i = 14;

    operand_b_i = 20;

    #10;

    operand_a_i = 10;

    operand_b_i = 9;

    #10;

    operand_a_i = 6;

    operand_b_i = 20;

    #10;

    operand_a_i = 18;

    operand_b_i = 5;

    #10;

    operand_a_i = 1;

    operand_b_i = 15;

    #10;

    operand_a_i = 20;

    operand_b_i = 11;

    #10;

    operand_a_i = 14;

    operand_b_i = 19;

    #10;

    operand_a_i = 9;

    operand_b_i = 16;

    #10;

    operand_a_i = 14;

    operand_b_i = 15;

    #10;

    operand_a_i = 8;

    operand_b_i = 3;

    #10;

    operand_a_i = 20;

    operand_b_i = 19;

    #10;

    operand_a_i = 20;

    operand_b_i = 17;

    #10;

    operand_a_i = 15;

    operand_b_i = 6;

    #10;

    operand_a_i = 13;

    operand_b_i = 14;

    #10;

    operand_a_i = 14;

    operand_b_i = 5;

    #10;

    operand_a_i = 3;

    operand_b_i = 11;

    #10;

    operand_a_i = 8;

    operand_b_i = 4;

    #10;

    operand_a_i = 19;

    operand_b_i = 14;

    #10;

    operand_a_i = 16;

    operand_b_i = 7;

    #10;

    operand_a_i = 9;

    operand_b_i = 11;

    #10;

    operand_a_i = 12;

    operand_b_i = 17;

    #10;

    operand_a_i = 8;

    operand_b_i = 17;

    #10;

    operand_a_i = 5;

    operand_b_i = 4;

    #10;

    operand_a_i = 19;

    operand_b_i = 16;

    #10;

    operand_a_i = 12;

    operand_b_i = 10;

    #10;

    operand_a_i = 13;

    operand_b_i = 14;

    #10;

    operand_a_i = 9;

    operand_b_i = 1;

    #10;

    operand_a_i = 8;

    operand_b_i = 5;

    #10;

    operand_a_i = 15;

    operand_b_i = 6;

    #10;

    operand_a_i = 2;

    operand_b_i = 15;

    #10;

    operand_a_i = 10;

    operand_b_i = 5;

    #10;

    operand_a_i = 1;

    operand_b_i = 5;

    #10;

    operand_a_i = 17;

    operand_b_i = 18;

    #10;

    operand_a_i = 2;

    operand_b_i = 9;

    #10;

    operand_a_i = 10;

    operand_b_i = 12;

    #10;

    operand_a_i = 14;

    operand_b_i = 10;

    #10;

    operand_a_i = 14;

    operand_b_i = 18;

    #10;

    operand_a_i = 11;

    operand_b_i = 4;

    #10;

    operand_a_i = 4;

    operand_b_i = 15;

    #10;

    operand_a_i = 10;

    operand_b_i = 18;

    #10;

    operand_a_i = 18;

    operand_b_i = 1;

    #10;

    operand_a_i = 3;

    operand_b_i = 18;

    #10;

    operand_a_i = 17;

    operand_b_i = 3;

    #10;

    operand_a_i = 5;

    operand_b_i = 16;

    #10;

    operand_a_i = 2;

    operand_b_i = 6;

    #10;

    operand_a_i = 15;

    operand_b_i = 18;

    #10;

    operand_a_i = 20;

    operand_b_i = 14;

    #10;

    operand_a_i = 8;

    operand_b_i = 1;

    #10;

    operand_a_i = 11;

    operand_b_i = 5;

    #10;

    operand_a_i = 7;

    operand_b_i = 3;

    #10;

    operand_a_i = 10;

    operand_b_i = 5;

    #10;

    operand_a_i = 5;

    operand_b_i = 4;

    #10;

    operand_a_i = 5;

    operand_b_i = 19;

    #10;

    operand_a_i = 3;

    operand_b_i = 20;

    #10;

    operand_a_i = 15;

    operand_b_i = 12;

    #10;

    operand_a_i = 9;

    operand_b_i = 15;

    #10;

    operand_a_i = 18;

    operand_b_i = 8;

    #10;

    operand_a_i = 3;

    operand_b_i = 14;

    #10;

    operand_a_i = 8;

    operand_b_i = 2;

    #10;

    operand_a_i = 10;

    operand_b_i = 20;

    #10;

    operand_a_i = 3;

    operand_b_i = 9;

    #10;

    operand_a_i = 5;

    operand_b_i = 15;

    #10;

    operand_a_i = 1;

    operand_b_i = 4;

    #10;

    operand_a_i = 2;

    operand_b_i = 3;

    #10;

    operand_a_i = 7;

    operand_b_i = 9;

    #10;

    operand_a_i = 3;

    operand_b_i = 19;

    #10;

    operand_a_i = 18;

    operand_b_i = 7;

    #10;

    operand_a_i = 13;

    operand_b_i = 6;

    #10;

    operand_a_i = 10;

    operand_b_i = 1;

    #10;

    operand_a_i = 9;

    operand_b_i = 1;

    #10;

    operand_a_i = 4;

    operand_b_i = 12;

    #10;

    operand_a_i = 2;

    operand_b_i = 20;

    #10;

    operand_a_i = 7;

    operand_b_i = 11;

    #10;

    operand_a_i = 10;

    operand_b_i = 4;

    #10;

    operand_a_i = 13;

    operand_b_i = 7;

    #10;

    operand_a_i = 20;

    operand_b_i = 3;

    #10;

    operand_a_i = 1;

    operand_b_i = 8;

    #10;

    operand_a_i = 18;

    operand_b_i = 4;

    #10;

    operand_a_i = 17;

    operand_b_i = 18;

    #10;

    operand_a_i = 7;

    operand_b_i = 5;

    #10;

    operand_a_i = 11;

    operand_b_i = 3;

    #10;

    operand_a_i = 15;

    operand_b_i = 9;

    #10;

    operand_a_i = 13;

    operand_b_i = 10;

    #10;

    operand_a_i = 11;

    operand_b_i = 16;

    #10;

    operand_a_i = 8;

    operand_b_i = 11;

    #10;

    operand_a_i = 4;

    operand_b_i = 3;

    #10;

    operand_a_i = 13;

    operand_b_i = 10;

    #10;

    operand_a_i = 10;

    operand_b_i = 11;

    #10;

    operand_a_i = 16;

    operand_b_i = 5;

    #10;

    operand_a_i = 12;

    operand_b_i = 3;

    #10;

    operand_a_i = 15;

    operand_b_i = 14;

    #10;

    operand_a_i = 8;

    operand_b_i = 19;

    #10;

    operand_a_i = 11;

    operand_b_i = 2;

    #10;

    operand_a_i = 2;

    operand_b_i = 6;

    #10;

    operand_a_i = 20;

    operand_b_i = 12;

    #10;

    operand_a_i = 3;

    operand_b_i = 12;

    #10;

    operand_a_i = 17;

    operand_b_i = 10;

    #10;

    operand_a_i = 14;

    operand_b_i = 19;

    #10;

    operand_a_i = 3;

    operand_b_i = 2;

    #10;

    operand_a_i = 10;

    operand_b_i = 7;

    #10;

    operand_a_i = 12;

    operand_b_i = 5;

    #10;

    operand_a_i = 2;

    operand_b_i = 18;

    #10;

    operand_a_i = 9;

    operand_b_i = 20;

    #10;

    operand_a_i = 12;

    operand_b_i = 9;

    #10;

    operand_a_i = 4;

    operand_b_i = 10;

    #10;

    operand_a_i = 18;

    operand_b_i = 3;

    #10;

    operand_a_i = 1;

    operand_b_i = 15;

    #10;

    operand_a_i = 10;

    operand_b_i = 11;

    #10;

    operand_a_i = 13;

    operand_b_i = 4;

    #10;

    operand_a_i = 15;

    operand_b_i = 11;

    #10;

    operand_a_i = 20;

    operand_b_i = 1;

    #10;

    operand_a_i = 2;

    operand_b_i = 9;

    #10;

    operand_a_i = 5;

    operand_b_i = 17;

    #10;

    operand_a_i = 15;

    operand_b_i = 12;

    #10;

    operand_a_i = 14;

    operand_b_i = 2;

    #10;

    operand_a_i = 3;

    operand_b_i = 7;

    #10;

    operand_a_i = 10;

    operand_b_i = 4;

    #10;

    operand_a_i = 4;

    operand_b_i = 2;

    #10;

    operand_a_i = 13;

    operand_b_i = 18;

    #10;

    operand_a_i = 14;

    operand_b_i = 3;

    #10;

    operand_a_i = 19;

    operand_b_i = 18;

    #10;

    operand_a_i = 1;

    operand_b_i = 7;

    #10;

    operand_a_i = 19;

    operand_b_i = 9;

    #10;

    operand_a_i = 2;

    operand_b_i = 15;

    #10;

    operand_a_i = 10;

    operand_b_i = 5;

    #10;

    operand_a_i = 14;

    operand_b_i = 19;

    #10;

    operand_a_i = 3;

    operand_b_i = 4;

    #10;

    operand_a_i = 15;

    operand_b_i = 12;

    #10;

    operand_a_i = 4;

    operand_b_i = 17;

    #10;

    operand_a_i = 1;

    operand_b_i = 15;

    #10;

    operand_a_i = 6;

    operand_b_i = 17;

    #10;

    operand_a_i = 9;

    operand_b_i = 20;

    #10;

    operand_a_i = 9;

    operand_b_i = 20;

    #10;

    operand_a_i = 1;

    operand_b_i = 15;

    #10;

    operand_a_i = 12;

    operand_b_i = 16;

    #10;

    operand_a_i = 9;

    operand_b_i = 13;

    #10;

    operand_a_i = 18;

    operand_b_i = 7;

    #10;

    operand_a_i = 11;

    operand_b_i = 2;

    #10;

    operand_a_i = 12;

    operand_b_i = 1;

    #10;

    operand_a_i = 19;

    operand_b_i = 13;

    #10;

    operand_a_i = 1;

    operand_b_i = 20;

    #10;

    operand_a_i = 5;

    operand_b_i = 17;

    #10;

    operand_a_i = 20;

    operand_b_i = 12;

    #10;

    operand_a_i = 15;

    operand_b_i = 11;

    #10;

    operand_a_i = 19;

    operand_b_i = 17;

    #10;

    operand_a_i = 1;

    operand_b_i = 14;

    #10;

    operand_a_i = 9;

    operand_b_i = 4;

    #10;

    operand_a_i = 17;

    operand_b_i = 4;

    #10;

    operand_a_i = 20;

    operand_b_i = 18;

    #10;

    operand_a_i = 6;

    operand_b_i = 4;

    #10;

    operand_a_i = 16;

    operand_b_i = 6;

    #10;

    operand_a_i = 14;

    operand_b_i = 16;

    #10;

    operand_a_i = 20;

    operand_b_i = 8;

    #10;

    operand_a_i = 9;

    operand_b_i = 8;

    #10;

    operand_a_i = 4;

    operand_b_i = 10;

    #10;

    operand_a_i = 17;

    operand_b_i = 9;

    #10;

    operand_a_i = 8;

    operand_b_i = 11;

    #10;

    operand_a_i = 7;

    operand_b_i = 12;

    #10;

    operand_a_i = 10;

    operand_b_i = 8;

    #10;

    operand_a_i = 9;

    operand_b_i = 15;

    #10;

    operand_a_i = 10;

    operand_b_i = 1;

    #10;

    operand_a_i = 7;

    operand_b_i = 8;

    #10;

    operand_a_i = 1;

    operand_b_i = 16;

    #10;

    operand_a_i = 7;

    operand_b_i = 17;

    #10;

    operand_a_i = 9;

    operand_b_i = 10;

    #10;

    operand_a_i = 7;

    operand_b_i = 14;

    #10;

    operand_a_i = 3;

    operand_b_i = 15;

    #10;

    operand_a_i = 11;

    operand_b_i = 10;

    #10;

    operand_a_i = 2;

    operand_b_i = 12;

    #10;

    operand_a_i = 18;

    operand_b_i = 6;

    #10;

    operand_a_i = 5;

    operand_b_i = 12;

    #10;

    operand_a_i = 20;

    operand_b_i = 11;

    #10;

    operand_a_i = 14;

    operand_b_i = 8;

    #10;

    operand_a_i = 17;

    operand_b_i = 2;

    #10;

    operand_a_i = 10;

    operand_b_i = 8;

    #10;

    operand_a_i = 7;

    operand_b_i = 16;

    #10;

    operand_a_i = 6;

    operand_b_i = 13;

    #10;

    operand_a_i = 18;

    operand_b_i = 13;

    #10;

    operand_a_i = 6;

    operand_b_i = 2;

    #10;

    operand_a_i = 3;

    operand_b_i = 1;

    #10;

    operand_a_i = 9;

    operand_b_i = 10;

    #10;

    operand_a_i = 12;

    operand_b_i = 6;

    #10;

    operand_a_i = 3;

    operand_b_i = 10;

    #10;

    operand_a_i = 2;

    operand_b_i = 3;

    #10;

    operand_a_i = 11;

    operand_b_i = 12;

    #10;

    operand_a_i = 16;

    operand_b_i = 8;

    #10;

    operand_a_i = 7;

    operand_b_i = 12;

    #10;

    operand_a_i = 8;

    operand_b_i = 13;

    #10;

    operand_a_i = 4;

    operand_b_i = 15;

    #10;

    operand_a_i = 5;

    operand_b_i = 13;

    #10;

    operand_a_i = 3;

    operand_b_i = 11;

    #10;

    operand_a_i = 14;

    operand_b_i = 13;

    #10;

    operand_a_i = 2;

    operand_b_i = 20;

    #10;

    operand_a_i = 9;

    operand_b_i = 5;

    #10;

    operand_a_i = 8;

    operand_b_i = 11;

    #10;

    operand_a_i = 1;

    operand_b_i = 14;

    #10;

    operand_a_i = 19;

    operand_b_i = 7;

    #10;

    operand_a_i = 16;

    operand_b_i = 19;

    #10;

    operand_a_i = 10;

    operand_b_i = 9;

    #10;

    operand_a_i = 16;

    operand_b_i = 7;

    #10;

    operand_a_i = 13;

    operand_b_i = 3;

    #10;

    operand_a_i = 11;

    operand_b_i = 10;

    #10;

    operand_a_i = 19;

    operand_b_i = 10;

    #10;

    operand_a_i = 5;

    operand_b_i = 4;

    #10;

    operand_a_i = 2;

    operand_b_i = 13;

    #10;

    operand_a_i = 10;

    operand_b_i = 18;

    #10;

    operand_a_i = 15;

    operand_b_i = 11;

    #10;

    operand_a_i = 3;

    operand_b_i = 10;

    #10;

    operand_a_i = 19;

    operand_b_i = 12;

    #10;

    operand_a_i = 10;

    operand_b_i = 13;

    #10;

    operand_a_i = 7;

    operand_b_i = 17;

    #10;

    operand_a_i = 12;

    operand_b_i = 15;

    #10;

    operand_a_i = 17;

    operand_b_i = 10;

    #10;

    operand_a_i = 7;

    operand_b_i = 5;

    #10;

    operand_a_i = 16;

    operand_b_i = 17;

    #10;

    operand_a_i = 15;

    operand_b_i = 2;

    #10;

    operand_a_i = 4;

    operand_b_i = 19;

    #10;

    operand_a_i = 13;

    operand_b_i = 2;

    #10;

    operand_a_i = 5;

    operand_b_i = 3;

    #10;

    operand_a_i = 1;

    operand_b_i = 13;

    #10;

    operand_a_i = 17;

    operand_b_i = 16;

    #10;

    operand_a_i = 4;

    operand_b_i = 11;

    #10;

    operand_a_i = 13;

    operand_b_i = 2;

    #10;

    operand_a_i = 7;

    operand_b_i = 12;

    #10;

    operand_a_i = 18;

    operand_b_i = 20;

    #10;

    operand_a_i = 11;

    operand_b_i = 14;

    #10;

    operand_a_i = 18;

    operand_b_i = 15;

    #10;

    operand_a_i = 3;

    operand_b_i = 17;

    #10;

    operand_a_i = 14;

    operand_b_i = 18;

    #10;

    operand_a_i = 4;

    operand_b_i = 6;

    #10;

    operand_a_i = 8;

    operand_b_i = 17;

    #10;

    operand_a_i = 12;

    operand_b_i = 10;

    #10;

    operand_a_i = 2;

    operand_b_i = 13;

    #10;

    operand_a_i = 14;

    operand_b_i = 8;

    #10;

    operand_a_i = 9;

    operand_b_i = 2;

    #10;

    operand_a_i = 5;

    operand_b_i = 11;

    #10;

    operand_a_i = 7;

    operand_b_i = 9;

    #10;

    operand_a_i = 17;

    operand_b_i = 20;

    #10;

    operand_a_i = 15;

    operand_b_i = 2;

    #10;

    operand_a_i = 16;

    operand_b_i = 9;

    #10;

    operand_a_i = 10;

    operand_b_i = 14;

    #10;

    operand_a_i = 1;

    operand_b_i = 5;

    #10;

    operand_a_i = 12;

    operand_b_i = 19;

    #10;

    operand_a_i = 11;

    operand_b_i = 2;

    #10;

    operand_a_i = 7;

    operand_b_i = 14;

    #10;

    operand_a_i = 9;

    operand_b_i = 16;

    #10;

    operand_a_i = 19;

    operand_b_i = 13;

    #10;

    operand_a_i = 10;

    operand_b_i = 12;

    #10;

    operand_a_i = 14;

    operand_b_i = 4;

    #10;

    operand_a_i = 2;

    operand_b_i = 6;

    #10;

    operand_a_i = 3;

    operand_b_i = 11;

    #10;

    operand_a_i = 4;

    operand_b_i = 20;

    #10;

    operand_a_i = 8;

    operand_b_i = 2;

    #10;

    operand_a_i = 14;

    operand_b_i = 15;

    #10;

    operand_a_i = 8;

    operand_b_i = 16;

    #10;

    operand_a_i = 11;

    operand_b_i = 5;

    #10;

    operand_a_i = 4;

    operand_b_i = 11;

    #10;

    operand_a_i = 9;

    operand_b_i = 19;

    #10;

    operand_a_i = 3;

    operand_b_i = 1;

    #10;

    operand_a_i = 14;

    operand_b_i = 6;

    #10;

    operand_a_i = 5;

    operand_b_i = 16;

    #10;

    operand_a_i = 15;

    operand_b_i = 9;

    #10;

    operand_a_i = 17;

    operand_b_i = 11;

    #10;

    operand_a_i = 10;

    operand_b_i = 20;

    #10;

    operand_a_i = 4;

    operand_b_i = 3;

    #10;

    operand_a_i = 14;

    operand_b_i = 4;

    #10;

    operand_a_i = 4;

    operand_b_i = 15;

    #10;

    operand_a_i = 12;

    operand_b_i = 2;

    #10;

    operand_a_i = 5;

    operand_b_i = 3;

    #10;

    operand_a_i = 5;

    operand_b_i = 17;

    #10;

    operand_a_i = 18;

    operand_b_i = 20;

    #10;

    operand_a_i = 15;

    operand_b_i = 14;

    #10;

    operand_a_i = 8;

    operand_b_i = 16;

    #10;

    operand_a_i = 13;

    operand_b_i = 8;

    #10;

    operand_a_i = 18;

    operand_b_i = 14;

    #10;

    operand_a_i = 5;

    operand_b_i = 15;

    #10;

    operand_a_i = 7;

    operand_b_i = 3;

    #10;

    operand_a_i = 10;

    operand_b_i = 1;

    #10;

    operand_a_i = 17;

    operand_b_i = 8;

    #10;

    operand_a_i = 7;

    operand_b_i = 10;

    #10;

    operand_a_i = 9;

    operand_b_i = 20;

    #10;

    operand_a_i = 16;

    operand_b_i = 4;

    #10;

    operand_a_i = 9;

    operand_b_i = 6;

    #10;

    operand_a_i = 6;

    operand_b_i = 14;

    #10;

    operand_a_i = 3;

    operand_b_i = 7;

    #10;

    operand_a_i = 4;

    operand_b_i = 9;

    #10;

    operand_a_i = 14;

    operand_b_i = 2;

    #10;

    operand_a_i = 13;

    operand_b_i = 10;

    #10;

    operand_a_i = 4;

    operand_b_i = 20;

    #10;

    operand_a_i = 12;

    operand_b_i = 15;

    #10;

    operand_a_i = 3;

    operand_b_i = 18;

    #10;

    operand_a_i = 12;

    operand_b_i = 16;

    #10;

    operand_a_i = 1;

    operand_b_i = 8;

    #10;

    operand_a_i = 8;

    operand_b_i = 12;

    #10;

    operand_a_i = 13;

    operand_b_i = 17;

    #10;

    operand_a_i = 20;

    operand_b_i = 15;

    #10;

    operand_a_i = 14;

    operand_b_i = 2;

    #10;

    operand_a_i = 17;

    operand_b_i = 6;

    #10;

    operand_a_i = 6;

    operand_b_i = 11;

    #10;

    operand_a_i = 18;

    operand_b_i = 4;

    #10;

    operand_a_i = 13;

    operand_b_i = 9;

    #10;

    operand_a_i = 7;

    operand_b_i = 6;

    #10;

    operand_a_i = 17;

    operand_b_i = 4;

    #10;

    operand_a_i = 3;

    operand_b_i = 12;

    #10;

    operand_a_i = 14;

    operand_b_i = 17;

    #10;

    operand_a_i = 13;

    operand_b_i = 4;

    #10;

    operand_a_i = 17;

    operand_b_i = 10;

    #10;

    operand_a_i = 10;

    operand_b_i = 3;

    #10;

    operand_a_i = 17;

    operand_b_i = 1;

    #10;

    operand_a_i = 13;

    operand_b_i = 8;

    #10;

    operand_a_i = 16;

    operand_b_i = 17;

    #10;

    operand_a_i = 7;

    operand_b_i = 5;

    #10;

    operand_a_i = 7;

    operand_b_i = 4;

    #10;

    operand_a_i = 7;

    operand_b_i = 13;

    #10;

    operand_a_i = 16;

    operand_b_i = 13;

    #10;

    operand_a_i = 16;

    operand_b_i = 19;

    #10;

    operand_a_i = 10;

    operand_b_i = 9;

    #10;

    operand_a_i = 9;

    operand_b_i = 19;

    #10;

    operand_a_i = 3;

    operand_b_i = 8;

    #10;

    operand_a_i = 15;

    operand_b_i = 5;

    #10;

    operand_a_i = 2;

    operand_b_i = 18;

    #10;

    operand_a_i = 3;

    operand_b_i = 10;

    #10;

    operand_a_i = 7;

    operand_b_i = 16;

    #10;

    operand_a_i = 6;

    operand_b_i = 20;

    #10;

    operand_a_i = 3;

    operand_b_i = 9;

    #10;

    operand_a_i = 19;

    operand_b_i = 5;

    #10;

    operand_a_i = 4;

    operand_b_i = 8;

    #10;

    operand_a_i = 8;

    operand_b_i = 10;

    #10;

    operand_a_i = 6;

    operand_b_i = 17;

    #10;

    operand_a_i = 7;

    operand_b_i = 14;

    #10;

    operand_a_i = 4;

    operand_b_i = 2;

    #10;

    operand_a_i = 1;

    operand_b_i = 3;

    #10;

    operand_a_i = 19;

    operand_b_i = 1;

    #10;

    operand_a_i = 15;

    operand_b_i = 20;

    #10;

    operand_a_i = 14;

    operand_b_i = 11;

    #10;

    operand_a_i = 6;

    operand_b_i = 9;

    #10;

    operand_a_i = 11;

    operand_b_i = 19;

    #10;

    operand_a_i = 19;

    operand_b_i = 13;

    #10;

    operand_a_i = 14;

    operand_b_i = 19;

    #10;

    operand_a_i = 19;

    operand_b_i = 1;

    #10;

    operand_a_i = 16;

    operand_b_i = 18;

    #10;

    operand_a_i = 18;

    operand_b_i = 10;

    #10;

    operand_a_i = 4;

    operand_b_i = 14;

    #10;

    operand_a_i = 11;

    operand_b_i = 17;

    #10;

    operand_a_i = 10;

    operand_b_i = 6;

    #10;

    operand_a_i = 14;

    operand_b_i = 6;

    #10;

    operand_a_i = 7;

    operand_b_i = 3;

    #10;

    operand_a_i = 6;

    operand_b_i = 3;

    #10;

    operand_a_i = 12;

    operand_b_i = 10;

    #10;

    operand_a_i = 1;

    operand_b_i = 14;

    #10;

    operand_a_i = 8;

    operand_b_i = 18;

    #10;

    operand_a_i = 10;

    operand_b_i = 14;

    #10;

    operand_a_i = 4;

    operand_b_i = 15;

    #10;

    operand_a_i = 17;

    operand_b_i = 13;

    #10;

    operand_a_i = 7;

    operand_b_i = 14;

    #10;

    operand_a_i = 5;

    operand_b_i = 19;

    #10;

    operand_a_i = 17;

    operand_b_i = 11;

    #10;

    operand_a_i = 1;

    operand_b_i = 19;

    #10;

    operand_a_i = 17;

    operand_b_i = 3;

    #10;

    operand_a_i = 9;

    operand_b_i = 5;

    #10;

    operand_a_i = 6;

    operand_b_i = 11;

    #10;

    operand_a_i = 7;

    operand_b_i = 4;

    #10;

    operand_a_i = 17;

    operand_b_i = 14;

    #10;

    operand_a_i = 19;

    operand_b_i = 11;

    #10;

    operand_a_i = 6;

    operand_b_i = 2;

    #10;

    operand_a_i = 13;

    operand_b_i = 17;

    #10;

    operand_a_i = 12;

    operand_b_i = 2;

    #10;

    operand_a_i = 20;

    operand_b_i = 16;

    #10;

    operand_a_i = 12;

    operand_b_i = 7;

    #10;

    operand_a_i = 14;

    operand_b_i = 8;

    #10;

    operand_a_i = 7;

    operand_b_i = 5;

    #10;

    operand_a_i = 19;

    operand_b_i = 9;

    #10;

    operand_a_i = 16;

    operand_b_i = 8;

    #10;

    operand_a_i = 4;

    operand_b_i = 14;

    #10;

    operand_a_i = 20;

    operand_b_i = 18;

    #10;

    operand_a_i = 18;

    operand_b_i = 14;

    #10;

    operand_a_i = 3;

    operand_b_i = 2;

    #10;

    operand_a_i = 18;

    operand_b_i = 20;

    #10;

    operand_a_i = 7;

    operand_b_i = 11;

    #10;

    operand_a_i = 17;

    operand_b_i = 3;

    #10;

    operand_a_i = 2;

    operand_b_i = 7;

    #10;

    operand_a_i = 4;

    operand_b_i = 12;

    #10;

    operand_a_i = 11;

    operand_b_i = 3;

    #10;

    operand_a_i = 13;

    operand_b_i = 10;

    #10;

    operand_a_i = 12;

    operand_b_i = 16;

    #10;

    operand_a_i = 13;

    operand_b_i = 3;

    #10;

    operand_a_i = 16;

    operand_b_i = 12;

    #10;

    operand_a_i = 6;

    operand_b_i = 9;

    #10;

    operand_a_i = 2;

    operand_b_i = 18;

    #10;

    operand_a_i = 16;

    operand_b_i = 6;

    #10;

    operand_a_i = 16;

    operand_b_i = 14;

    #10;

    operand_a_i = 14;

    operand_b_i = 3;

    #10;

    operand_a_i = 10;

    operand_b_i = 3;

    #10;

    operand_a_i = 2;

    operand_b_i = 12;

    #10;

    operand_a_i = 8;

    operand_b_i = 14;

    #10;

    operand_a_i = 16;

    operand_b_i = 1;

    #10;

    operand_a_i = 5;

    operand_b_i = 12;

    #10;

    operand_a_i = 19;

    operand_b_i = 8;

    #10;

    operand_a_i = 14;

    operand_b_i = 16;

    #10;

    operand_a_i = 12;

    operand_b_i = 7;

    #10;

    operand_a_i = 11;

    operand_b_i = 10;

    #10;

    operand_a_i = 9;

    operand_b_i = 8;

    #10;

    operand_a_i = 15;

    operand_b_i = 1;

    #10;

    operand_a_i = 19;

    operand_b_i = 4;

    #10;

    operand_a_i = 18;

    operand_b_i = 16;

    #10;

    operand_a_i = 12;

    operand_b_i = 4;

    #10;

    operand_a_i = 17;

    operand_b_i = 8;

    #10;

    operand_a_i = 11;

    operand_b_i = 6;

    #10;

    operand_a_i = 18;

    operand_b_i = 10;

    #10;

    operand_a_i = 19;

    operand_b_i = 12;

    #10;

    operand_a_i = 11;

    operand_b_i = 18;

    #10;

    operand_a_i = 5;

    operand_b_i = 7;

    #10;

    operand_a_i = 11;

    operand_b_i = 8;

    #10;

    operand_a_i = 14;

    operand_b_i = 8;

    #10;

    operand_a_i = 2;

    operand_b_i = 4;

    #10;

    operand_a_i = 10;

    operand_b_i = 5;

    #10;

    operand_a_i = 2;

    operand_b_i = 17;

    #10;

    operand_a_i = 12;

    operand_b_i = 15;

    #10;

    operand_a_i = 15;

    operand_b_i = 10;

    #10;

    operand_a_i = 15;

    operand_b_i = 19;

    #10;

    operand_a_i = 7;

    operand_b_i = 12;

    #10;

    operand_a_i = 5;

    operand_b_i = 16;

    #10;

    operand_a_i = 15;

    operand_b_i = 10;

    #10;

    operand_a_i = 15;

    operand_b_i = 7;

    #10;

    operand_a_i = 10;

    operand_b_i = 8;

    #10;

    operand_a_i = 15;

    operand_b_i = 1;

    #10;

    operand_a_i = 18;

    operand_b_i = 6;

    #10;

    operand_a_i = 4;

    operand_b_i = 18;

    #10;

    operand_a_i = 7;

    operand_b_i = 3;

    #10;

    operand_a_i = 10;

    operand_b_i = 6;

    #10;

    operand_a_i = 8;

    operand_b_i = 14;

    #10;

    operand_a_i = 7;

    operand_b_i = 1;

    #10;

    operand_a_i = 8;

    operand_b_i = 1;

    #10;

    operand_a_i = 17;

    operand_b_i = 5;

    #10;

    operand_a_i = 6;

    operand_b_i = 2;

    #10;

    operand_a_i = 7;

    operand_b_i = 14;

    #10;

    operand_a_i = 15;

    operand_b_i = 6;

    #10;

    operand_a_i = 20;

    operand_b_i = 16;

    #10;

    operand_a_i = 4;

    operand_b_i = 8;

    #10;

    operand_a_i = 3;

    operand_b_i = 7;

    #10;

    operand_a_i = 14;

    operand_b_i = 8;

    #10;

    operand_a_i = 2;

    operand_b_i = 15;

    #10;

    operand_a_i = 6;

    operand_b_i = 9;

    #10;

    operand_a_i = 4;

    operand_b_i = 1;

    #10;

    operand_a_i = 5;

    operand_b_i = 8;

    #10;

    operand_a_i = 9;

    operand_b_i = 17;

    #10;

    operand_a_i = 20;

    operand_b_i = 1;

    #10;

    operand_a_i = 8;

    operand_b_i = 1;

    #10;

    operand_a_i = 19;

    operand_b_i = 18;

    #10;

    operand_a_i = 7;

    operand_b_i = 18;

    #10;

    operand_a_i = 8;

    operand_b_i = 11;

    #10;

    operand_a_i = 9;

    operand_b_i = 6;

    #10;

    operand_a_i = 1;

    operand_b_i = 20;

    #10;

    operand_a_i = 12;

    operand_b_i = 3;

    #10;

    operand_a_i = 5;

    operand_b_i = 6;

    #10;

    operand_a_i = 6;

    operand_b_i = 9;

    #10;

    operand_a_i = 16;

    operand_b_i = 18;

    #10;

    operand_a_i = 13;

    operand_b_i = 1;

    #10;

    operand_a_i = 11;

    operand_b_i = 13;

    #10;

    operand_a_i = 18;

    operand_b_i = 2;

    #10;

    operand_a_i = 11;

    operand_b_i = 19;

    #10;

    operand_a_i = 7;

    operand_b_i = 11;

    #10;

    operand_a_i = 20;

    operand_b_i = 5;

    #10;

    operand_a_i = 2;

    operand_b_i = 7;

    #10;

    operand_a_i = 17;

    operand_b_i = 8;

    #10;

    operand_a_i = 20;

    operand_b_i = 12;

    #10;

    operand_a_i = 19;

    operand_b_i = 3;

    #10;

    operand_a_i = 2;

    operand_b_i = 11;

    #10;

    operand_a_i = 18;

    operand_b_i = 20;

    #10;

    operand_a_i = 3;

    operand_b_i = 5;

    #10;

    operand_a_i = 19;

    operand_b_i = 1;

    #10;

    operand_a_i = 5;

    operand_b_i = 18;

    #10;

    operand_a_i = 5;

    operand_b_i = 13;

    #10;

    operand_a_i = 3;

    operand_b_i = 17;

    #10;

    operand_a_i = 9;

    operand_b_i = 16;

    #10;

    operand_a_i = 6;

    operand_b_i = 16;

    #10;

    operand_a_i = 11;

    operand_b_i = 9;

    #10;

    operand_a_i = 2;

    operand_b_i = 11;

    #10;

    operand_a_i = 13;

    operand_b_i = 18;

    #10;

    operand_a_i = 20;

    operand_b_i = 17;

    #10;

    operand_a_i = 7;

    operand_b_i = 14;

    #10;

    operand_a_i = 4;

    operand_b_i = 6;

    #10;

    operand_a_i = 18;

    operand_b_i = 19;

    #10;

    operand_a_i = 20;

    operand_b_i = 17;

    #10;

    operand_a_i = 19;

    operand_b_i = 7;

    #10;

    operand_a_i = 6;

    operand_b_i = 11;

    #10;

    operand_a_i = 17;

    operand_b_i = 10;

    #10;

    operand_a_i = 20;

    operand_b_i = 12;

    #10;

    operand_a_i = 7;

    operand_b_i = 10;

    #10;

    operand_a_i = 20;

    operand_b_i = 15;

    #10;

    operand_a_i = 3;

    operand_b_i = 14;

    #10;

    operand_a_i = 14;

    operand_b_i = 3;

    #10;

    operand_a_i = 6;

    operand_b_i = 8;

    #10;

    operand_a_i = 13;

    operand_b_i = 11;

    #10;

    operand_a_i = 14;

    operand_b_i = 4;

    #10;

    operand_a_i = 1;

    operand_b_i = 2;

    #10;

    operand_a_i = 2;

    operand_b_i = 7;

    #10;

    operand_a_i = 6;

    operand_b_i = 3;

    #10;

    operand_a_i = 6;

    operand_b_i = 13;

    #10;

    operand_a_i = 4;

    operand_b_i = 12;

    #10;

    operand_a_i = 2;

    operand_b_i = 15;

    #10;

    operand_a_i = 1;

    operand_b_i = 17;

    #10;

    operand_a_i = 14;

    operand_b_i = 8;

    #10;

    operand_a_i = 4;

    operand_b_i = 12;

    #10;

    operand_a_i = 11;

    operand_b_i = 14;

    #10;

    operand_a_i = 4;

    operand_b_i = 18;

    #10;

    operand_a_i = 20;

    operand_b_i = 6;

    #10;

    operand_a_i = 1;

    operand_b_i = 9;

    #10;

    operand_a_i = 12;

    operand_b_i = 2;

    #10;

    operand_a_i = 14;

    operand_b_i = 5;

    #10;

    operand_a_i = 10;

    operand_b_i = 7;

    #10;

    operand_a_i = 9;

    operand_b_i = 17;

    #10;

    operand_a_i = 12;

    operand_b_i = 9;

    #10;

    operand_a_i = 9;

    operand_b_i = 13;

    #10;

    operand_a_i = 3;

    operand_b_i = 1;

    #10;

    operand_a_i = 4;

    operand_b_i = 20;

    #10;

    operand_a_i = 17;

    operand_b_i = 11;

    #10;

    operand_a_i = 17;

    operand_b_i = 2;

    #10;

    operand_a_i = 2;

    operand_b_i = 7;

    #10;

    operand_a_i = 13;

    operand_b_i = 17;

    #10;

    operand_a_i = 16;

    operand_b_i = 12;

    #10;

    operand_a_i = 10;

    operand_b_i = 16;

    #10;

    operand_a_i = 2;

    operand_b_i = 5;

    #10;

    operand_a_i = 19;

    operand_b_i = 10;

    #10;

    operand_a_i = 1;

    operand_b_i = 14;

    #10;

    operand_a_i = 6;

    operand_b_i = 19;

    #10;

    operand_a_i = 1;

    operand_b_i = 15;

    #10;

    operand_a_i = 4;

    operand_b_i = 15;

    #10;

    operand_a_i = 3;

    operand_b_i = 17;

    #10;

    operand_a_i = 15;

    operand_b_i = 12;

    #10;

    operand_a_i = 20;

    operand_b_i = 7;

    #10;

    operand_a_i = 10;

    operand_b_i = 4;

    #10;

    operand_a_i = 6;

    operand_b_i = 13;

    #10;

    operand_a_i = 12;

    operand_b_i = 6;

    #10;

    operand_a_i = 20;

    operand_b_i = 4;

    #10;

    operand_a_i = 3;

    operand_b_i = 11;

    #10;

    operand_a_i = 5;

    operand_b_i = 18;

    #10;

    operand_a_i = 6;

    operand_b_i = 16;

    #10;

    operand_a_i = 11;

    operand_b_i = 6;

    #10;

    operand_a_i = 19;

    operand_b_i = 17;

    #10;

    operand_a_i = 15;

    operand_b_i = 12;

    #10;

    operand_a_i = 17;

    operand_b_i = 12;

    #10;

    operand_a_i = 13;

    operand_b_i = 7;

    #10;

    operand_a_i = 5;

    operand_b_i = 17;

    #10;

    operand_a_i = 3;

    operand_b_i = 9;

    #10;

    operand_a_i = 3;

    operand_b_i = 14;

    #10;

    operand_a_i = 1;

    operand_b_i = 16;

    #10;

    operand_a_i = 12;

    operand_b_i = 14;

    #10;

    operand_a_i = 8;

    operand_b_i = 11;

    #10;

    operand_a_i = 11;

    operand_b_i = 3;

    #10;

    operand_a_i = 6;

    operand_b_i = 14;

    #10;

    operand_a_i = 4;

    operand_b_i = 5;

    #10;

    operand_a_i = 11;

    operand_b_i = 13;

    #10;

    operand_a_i = 12;

    operand_b_i = 6;

    #10;

    operand_a_i = 6;

    operand_b_i = 20;

    #10;

    operand_a_i = 14;

    operand_b_i = 19;

    #10;

    operand_a_i = 17;

    operand_b_i = 5;

    #10;

    operand_a_i = 15;

    operand_b_i = 4;

    #10;

    operand_a_i = 5;

    operand_b_i = 10;

    #10;

    operand_a_i = 20;

    operand_b_i = 9;

    #10;

    operand_a_i = 17;

    operand_b_i = 15;

    #10;

    operand_a_i = 11;

    operand_b_i = 16;

    #10;

    operand_a_i = 11;

    operand_b_i = 1;

    #10;

    operand_a_i = 3;

    operand_b_i = 18;

    #10;

    operand_a_i = 8;

    operand_b_i = 7;

    #10;

    operand_a_i = 9;

    operand_b_i = 12;

    #10;

    operand_a_i = 3;

    operand_b_i = 7;

    #10;

    operand_a_i = 3;

    operand_b_i = 8;

    #10;

    operand_a_i = 5;

    operand_b_i = 6;

    #10;

    operand_a_i = 19;

    operand_b_i = 5;

    #10;

    operand_a_i = 9;

    operand_b_i = 13;

    #10;

    operand_a_i = 5;

    operand_b_i = 4;

    #10;

    operand_a_i = 1;

    operand_b_i = 7;

    #10;

    operand_a_i = 18;

    operand_b_i = 16;

    #10;

    operand_a_i = 4;

    operand_b_i = 1;

    #10;

    operand_a_i = 2;

    operand_b_i = 15;

    #10;

    operand_a_i = 12;

    operand_b_i = 15;

    #10;

    operand_a_i = 2;

    operand_b_i = 13;

    #10;

    operand_a_i = 14;

    operand_b_i = 2;

    #10;

    operand_a_i = 19;

    operand_b_i = 1;

    #10;

    operand_a_i = 13;

    operand_b_i = 19;

    #10;

    operand_a_i = 6;

    operand_b_i = 9;

    #10;

    operand_a_i = 20;

    operand_b_i = 9;

    #10;

    operand_a_i = 11;

    operand_b_i = 6;

    #10;

    operand_a_i = 12;

    operand_b_i = 7;

    #10;

    operand_a_i = 10;

    operand_b_i = 20;

    #10;

    operand_a_i = 5;

    operand_b_i = 11;

    #10;

    operand_a_i = 15;

    operand_b_i = 2;

    #10;

    operand_a_i = 6;

    operand_b_i = 2;

    #10;

    operand_a_i = 15;

    operand_b_i = 16;

    #10;

    operand_a_i = 14;

    operand_b_i = 7;

    #10;

    operand_a_i = 12;

    operand_b_i = 3;

    #10;

    operand_a_i = 2;

    operand_b_i = 6;

    #10;

    operand_a_i = 1;

    operand_b_i = 14;

    #10;

    operand_a_i = 12;

    operand_b_i = 13;

    #10;

    operand_a_i = 16;

    operand_b_i = 2;

    #10;

    operand_a_i = 7;

    operand_b_i = 1;

    #10;

    operand_a_i = 3;

    operand_b_i = 6;

    #10;

    operand_a_i = 1;

    operand_b_i = 5;

    #10;

    operand_a_i = 16;

    operand_b_i = 10;

    #10;

    operand_a_i = 10;

    operand_b_i = 5;

    #10;

    operand_a_i = 7;

    operand_b_i = 15;

    #10;

    operand_a_i = 5;

    operand_b_i = 11;

    #10;

    operand_a_i = 10;

    operand_b_i = 4;

    #10;

    operand_a_i = 20;

    operand_b_i = 19;

    #10;

    operand_a_i = 8;

    operand_b_i = 15;

    #10;

    operand_a_i = 8;

    operand_b_i = 5;

    #10;

    operand_a_i = 14;

    operand_b_i = 3;

    #10;

    operand_a_i = 15;

    operand_b_i = 9;

    #10;

    operand_a_i = 12;

    operand_b_i = 18;

    #10;

    operand_a_i = 5;

    operand_b_i = 19;

    #10;

    operand_a_i = 19;

    operand_b_i = 18;

    #10;

    operand_a_i = 20;

    operand_b_i = 11;

    #10;

    operand_a_i = 12;

    operand_b_i = 19;

    #10;

    operand_a_i = 17;

    operand_b_i = 11;

    #10;

    operand_a_i = 17;

    operand_b_i = 16;

    #10;

    operand_a_i = 9;

    operand_b_i = 1;

    #10;

    operand_a_i = 3;

    operand_b_i = 6;

    #10;

    operand_a_i = 8;

    operand_b_i = 7;

    #10;

    operand_a_i = 11;

    operand_b_i = 13;

    #10;

    operand_a_i = 14;

    operand_b_i = 11;

    #10;

    operand_a_i = 6;

    operand_b_i = 16;

    #10;

    operand_a_i = 18;

    operand_b_i = 14;

    #10;

    operand_a_i = 20;

    operand_b_i = 2;

    #10;

    operand_a_i = 2;

    operand_b_i = 16;

    #10;

    operand_a_i = 7;

    operand_b_i = 13;

    #10;

    operand_a_i = 7;

    operand_b_i = 17;

    #10;

    operand_a_i = 15;

    operand_b_i = 12;

    #10;

    operand_a_i = 9;

    operand_b_i = 1;

    #10;

    operand_a_i = 18;

    operand_b_i = 15;

    #10;

    operand_a_i = 14;

    operand_b_i = 5;

    #10;

    operand_a_i = 4;

    operand_b_i = 3;

    #10;

    operand_a_i = 7;

    operand_b_i = 13;

    #10;

    operand_a_i = 10;

    operand_b_i = 1;

    #10;

    operand_a_i = 7;

    operand_b_i = 13;

    #10;

    operand_a_i = 6;

    operand_b_i = 1;

    #10;

    operand_a_i = 20;

    operand_b_i = 14;

    #10;

    operand_a_i = 14;

    operand_b_i = 13;

    #10;

    operand_a_i = 1;

    operand_b_i = 6;

    #10;

    operand_a_i = 8;

    operand_b_i = 6;

    #10;

    operand_a_i = 14;

    operand_b_i = 16;

    #10;

    operand_a_i = 14;

    operand_b_i = 20;

    #10;

    operand_a_i = 1;

    operand_b_i = 3;

    #10;

    operand_a_i = 19;

    operand_b_i = 20;

    #10;

    operand_a_i = 5;

    operand_b_i = 3;

    #10;

    operand_a_i = 12;

    operand_b_i = 18;

    #10;

    operand_a_i = 12;

    operand_b_i = 11;

    #10;

    operand_a_i = 12;

    operand_b_i = 18;

    #10;

    operand_a_i = 17;

    operand_b_i = 8;

    #10;

    operand_a_i = 15;

    operand_b_i = 7;

    #10;

    operand_a_i = 9;

    operand_b_i = 20;

    #10;

    operand_a_i = 15;

    operand_b_i = 12;

    #10;

    operand_a_i = 19;

    operand_b_i = 13;

    #10;

    operand_a_i = 2;

    operand_b_i = 6;

    #10;

    operand_a_i = 1;

    operand_b_i = 20;

    #10;

    operand_a_i = 20;

    operand_b_i = 1;

    #10;

    operand_a_i = 13;

    operand_b_i = 17;

    #10;

    operand_a_i = 6;

    operand_b_i = 4;

    #10;

    operand_a_i = 14;

    operand_b_i = 15;

    #10;

    operand_a_i = 20;

    operand_b_i = 15;

    #10;

    operand_a_i = 3;

    operand_b_i = 10;

    #10;

    operand_a_i = 20;

    operand_b_i = 6;

    #10;

    operand_a_i = 7;

    operand_b_i = 2;

    #10;

    operand_a_i = 2;

    operand_b_i = 11;

    #10;

    operand_a_i = 5;

    operand_b_i = 1;

    #10;

    operand_a_i = 12;

    operand_b_i = 8;

    #10;

    operand_a_i = 20;

    operand_b_i = 5;

    #10;

    operand_a_i = 18;

    operand_b_i = 17;

    #10;

    operand_a_i = 10;

    operand_b_i = 1;

    #10;

    operand_a_i = 20;

    operand_b_i = 3;

    #10;

    operand_a_i = 2;

    operand_b_i = 6;

    #10;

    operand_a_i = 20;

    operand_b_i = 9;

    #10;

    operand_a_i = 15;

    operand_b_i = 8;

    #10;

    operand_a_i = 7;

    operand_b_i = 13;

    #10;

    operand_a_i = 18;

    operand_b_i = 14;

    #10;

    operand_a_i = 12;

    operand_b_i = 13;

    #10;

    operand_a_i = 1;

    operand_b_i = 12;

    #10;

    operand_a_i = 5;

    operand_b_i = 6;

    #10;

    operand_a_i = 5;

    operand_b_i = 11;

    #10;

    operand_a_i = 9;

    operand_b_i = 11;

    #10;

    operand_a_i = 18;

    operand_b_i = 12;

    #10;

    operand_a_i = 13;

    operand_b_i = 19;

    #10;

    operand_a_i = 3;

    operand_b_i = 4;

    #10;

    operand_a_i = 2;

    operand_b_i = 10;

    #10;

    operand_a_i = 8;

    operand_b_i = 2;

    #10;

    operand_a_i = 2;

    operand_b_i = 16;

    #10;

    operand_a_i = 8;

    operand_b_i = 1;

    #10;

    operand_a_i = 13;

    operand_b_i = 6;

    #10;

    operand_a_i = 14;

    operand_b_i = 19;

    #10;

    operand_a_i = 1;

    operand_b_i = 4;

    #10;

    operand_a_i = 8;

    operand_b_i = 10;

    #10;

    operand_a_i = 6;

    operand_b_i = 5;

    #10;

    operand_a_i = 8;

    operand_b_i = 18;

    #10;

    operand_a_i = 3;

    operand_b_i = 18;

    #10;

    operand_a_i = 11;

    operand_b_i = 9;

    #10;

    operand_a_i = 1;

    operand_b_i = 4;

    #10;

    operand_a_i = 18;

    operand_b_i = 5;

    #10;

    operand_a_i = 20;

    operand_b_i = 19;

    #10;

    operand_a_i = 20;

    operand_b_i = 6;

    #10;

    operand_a_i = 8;

    operand_b_i = 17;

    #10;

    operand_a_i = 11;

    operand_b_i = 16;

    #10;

    operand_a_i = 1;

    operand_b_i = 16;

    #10;

    operand_a_i = 18;

    operand_b_i = 7;

    #10;

    operand_a_i = 5;

    operand_b_i = 18;

    #10;

    operand_a_i = 11;

    operand_b_i = 18;

    #10;

    operand_a_i = 3;

    operand_b_i = 18;

    #10;

    operand_a_i = 18;

    operand_b_i = 1;

    #10;

    operand_a_i = 13;

    operand_b_i = 6;

    #10;

    operand_a_i = 10;

    operand_b_i = 18;

    #10;

    operand_a_i = 16;

    operand_b_i = 19;

    #10;

    operand_a_i = 18;

    operand_b_i = 12;

    #10;

    operand_a_i = 2;

    operand_b_i = 3;

    #10;

    operand_a_i = 8;

    operand_b_i = 16;

    #10;

    operand_a_i = 7;

    operand_b_i = 12;

    #10;

    operand_a_i = 16;

    operand_b_i = 19;

    #10;

    operand_a_i = 5;

    operand_b_i = 6;

    #10;

    operand_a_i = 9;

    operand_b_i = 12;

    #10;

    operand_a_i = 3;

    operand_b_i = 15;

    #10;

    operand_a_i = 3;

    operand_b_i = 2;

    #10;

    operand_a_i = 5;

    operand_b_i = 19;

    #10;

    operand_a_i = 2;

    operand_b_i = 20;

    #10;

    operand_a_i = 8;

    operand_b_i = 2;

    #10;

    operand_a_i = 16;

    operand_b_i = 2;

    #10;

    operand_a_i = 3;

    operand_b_i = 7;

    #10;

    operand_a_i = 4;

    operand_b_i = 14;

    #10;

    operand_a_i = 2;

    operand_b_i = 17;

    #10;

    operand_a_i = 6;

    operand_b_i = 17;

    #10;

    operand_a_i = 1;

    operand_b_i = 8;

    #10;

    operand_a_i = 13;

    operand_b_i = 14;

    #10;

    operand_a_i = 20;

    operand_b_i = 7;

    #10;

    operand_a_i = 9;

    operand_b_i = 16;

    #10;

    operand_a_i = 11;

    operand_b_i = 10;

    #10;

    operand_a_i = 18;

    operand_b_i = 12;

    #10;

    operand_a_i = 13;

    operand_b_i = 16;

    #10;

    operand_a_i = 6;

    operand_b_i = 19;

    #10;

    operand_a_i = 15;

    operand_b_i = 20;

    #10;

    operand_a_i = 3;

    operand_b_i = 10;

    #10;

    operand_a_i = 10;

    operand_b_i = 5;

    #10;

    operand_a_i = 12;

    operand_b_i = 10;

    #10;

    operand_a_i = 8;

    operand_b_i = 1;

    #10;

    operand_a_i = 11;

    operand_b_i = 14;

    #10;

    operand_a_i = 10;

    operand_b_i = 6;

    #10;

    operand_a_i = 18;

    operand_b_i = 14;

    #10;

    operand_a_i = 17;

    operand_b_i = 10;

    #10;

    operand_a_i = 11;

    operand_b_i = 2;

    #10;

    operand_a_i = 7;

    operand_b_i = 4;

    #10;

    operand_a_i = 10;

    operand_b_i = 18;

    #10;

    operand_a_i = 1;

    operand_b_i = 20;

    #10;

    operand_a_i = 5;

    operand_b_i = 7;

    #10;

    operand_a_i = 9;

    operand_b_i = 11;

    #10;

    operand_a_i = 15;

    operand_b_i = 5;

    #10;

    operand_a_i = 14;

    operand_b_i = 6;

    #10;

    operand_a_i = 4;

    operand_b_i = 20;

    #10;

    operand_a_i = 18;

    operand_b_i = 5;

    #10;

    operand_a_i = 18;

    operand_b_i = 11;

    #10;

    operand_a_i = 16;

    operand_b_i = 12;

    #10;

    operand_a_i = 19;

    operand_b_i = 18;

    #10;

    operand_a_i = 4;

    operand_b_i = 1;

    #10;

    operand_a_i = 12;

    operand_b_i = 9;

    #10;

    operand_a_i = 9;

    operand_b_i = 8;

    #10;

    operand_a_i = 2;

    operand_b_i = 1;

    #10;

    operand_a_i = 2;

    operand_b_i = 9;

    #10;

    operand_a_i = 9;

    operand_b_i = 10;

    #10;

    operand_a_i = 15;

    operand_b_i = 4;

    #10;

    operand_a_i = 4;

    operand_b_i = 2;

    #10;

    operand_a_i = 18;

    operand_b_i = 12;

    #10;

    operand_a_i = 15;

    operand_b_i = 20;

    #10;

    operand_a_i = 12;

    operand_b_i = 10;

    #10;

    operand_a_i = 8;

    operand_b_i = 9;

    #10;

    operand_a_i = 6;

    operand_b_i = 12;

    #10;

    operand_a_i = 13;

    operand_b_i = 20;

    #10;

    operand_a_i = 12;

    operand_b_i = 13;

    #10;

    operand_a_i = 15;

    operand_b_i = 9;

    #10;

    operand_a_i = 9;

    operand_b_i = 17;

    #10;

    operand_a_i = 13;

    operand_b_i = 5;

    #10;

    operand_a_i = 7;

    operand_b_i = 3;

    #10;

    operand_a_i = 4;

    operand_b_i = 12;

    #10;

    operand_a_i = 7;

    operand_b_i = 16;

    #10;

    operand_a_i = 1;

    operand_b_i = 13;

    #10;

    operand_a_i = 6;

    operand_b_i = 8;

    #10;

    operand_a_i = 17;

    operand_b_i = 13;

    #10;

    operand_a_i = 7;

    operand_b_i = 14;

    #10;

    operand_a_i = 16;

    operand_b_i = 1;

    #10;

    operand_a_i = 9;

    operand_b_i = 4;

    #10;

    operand_a_i = 11;

    operand_b_i = 5;

    #10;

    operand_a_i = 6;

    operand_b_i = 13;

    #10;

    operand_a_i = 19;

    operand_b_i = 18;

    #10;

    operand_a_i = 20;

    operand_b_i = 5;

    #10;

    operand_a_i = 12;

    operand_b_i = 9;

    #10;

    operand_a_i = 15;

    operand_b_i = 20;

    #10;

    operand_a_i = 18;

    operand_b_i = 13;

    #10;

    operand_a_i = 18;

    operand_b_i = 15;

    #10;

    operand_a_i = 7;

    operand_b_i = 10;

    #10;

    operand_a_i = 13;

    operand_b_i = 14;

    #10;

    operand_a_i = 6;

    operand_b_i = 11;

    #10;

    operand_a_i = 1;

    operand_b_i = 6;

    #10;

    operand_a_i = 4;

    operand_b_i = 9;

    #10;

    operand_a_i = 8;

    operand_b_i = 6;

    #10;

    operand_a_i = 8;

    operand_b_i = 17;

    #10;

    operand_a_i = 15;

    operand_b_i = 8;

    #10;

    operand_a_i = 12;

    operand_b_i = 19;

    #10;

    operand_a_i = 6;

    operand_b_i = 14;

    #10;

    operand_a_i = 12;

    operand_b_i = 16;

    #10;

    operand_a_i = 2;

    operand_b_i = 20;

    #10;

    operand_a_i = 5;

    operand_b_i = 11;

    #10;

    operand_a_i = 12;

    operand_b_i = 7;

    #10;

    operand_a_i = 3;

    operand_b_i = 10;

    #10;

    operand_a_i = 12;

    operand_b_i = 2;

    #10;

    operand_a_i = 12;

    operand_b_i = 13;

    #10;

    operand_a_i = 3;

    operand_b_i = 19;

    #10;

    operand_a_i = 14;

    operand_b_i = 6;

    #10;

    operand_a_i = 6;

    operand_b_i = 14;

    #10;

    operand_a_i = 10;

    operand_b_i = 14;

    #10;

    operand_a_i = 15;

    operand_b_i = 6;

    #10;

    operand_a_i = 18;

    operand_b_i = 4;

    #10;

    operand_a_i = 18;

    operand_b_i = 20;

    #10;

    operand_a_i = 15;

    operand_b_i = 9;

    #10;

    operand_a_i = 9;

    operand_b_i = 17;

    #10;

    operand_a_i = 3;

    operand_b_i = 5;

    #10;

    operand_a_i = 4;

    operand_b_i = 19;

    #10;

    operand_a_i = 20;

    operand_b_i = 19;

    #10;

    operand_a_i = 1;

    operand_b_i = 9;

    #10;

    operand_a_i = 1;

    operand_b_i = 8;

    #10;

    operand_a_i = 6;

    operand_b_i = 12;

    #10;

    operand_a_i = 13;

    operand_b_i = 1;

    #10;

    operand_a_i = 13;

    operand_b_i = 5;

    #10;

    operand_a_i = 6;

    operand_b_i = 1;

    #10;

    operand_a_i = 14;

    operand_b_i = 20;

    #10;

    operand_a_i = 1;

    operand_b_i = 7;

    #10;

    operand_a_i = 5;

    operand_b_i = 1;

    #10;

    operand_a_i = 10;

    operand_b_i = 17;

    #10;

    operand_a_i = 15;

    operand_b_i = 5;

    #10;

    operand_a_i = 12;

    operand_b_i = 1;

    #10;

    operand_a_i = 2;

    operand_b_i = 3;

    #10;

    operand_a_i = 11;

    operand_b_i = 5;

    #10;

    operand_a_i = 1;

    operand_b_i = 12;

    #10;

    operand_a_i = 7;

    operand_b_i = 9;

    #10;

    operand_a_i = 12;

    operand_b_i = 13;

    #10;

    operand_a_i = 11;

    operand_b_i = 12;

    #10;

    operand_a_i = 1;

    operand_b_i = 6;

    #10;

    operand_a_i = 6;

    operand_b_i = 2;

    #10;

    operand_a_i = 13;

    operand_b_i = 19;

    #10;

    operand_a_i = 11;

    operand_b_i = 17;

    #10;

    operand_a_i = 17;

    operand_b_i = 5;

    #10;

    operand_a_i = 16;

    operand_b_i = 17;

    #10;

    operand_a_i = 14;

    operand_b_i = 6;

    #10;

    operand_a_i = 12;

    operand_b_i = 13;

    #10;

    operand_a_i = 8;

    operand_b_i = 7;

    #10;

    operand_a_i = 12;

    operand_b_i = 17;

    #10;

    operand_a_i = 2;

    operand_b_i = 4;

    #10;

    operand_a_i = 13;

    operand_b_i = 8;

    #10;

    operand_a_i = 10;

    operand_b_i = 16;

    #10;

    operand_a_i = 15;

    operand_b_i = 1;

    #10;

    operand_a_i = 19;

    operand_b_i = 12;

    #10;

    operand_a_i = 15;

    operand_b_i = 7;

    #10;

    operand_a_i = 5;

    operand_b_i = 12;

    #10;

    operand_a_i = 16;

    operand_b_i = 19;

    #10;

    operand_a_i = 6;

    operand_b_i = 8;

    #10;

    operand_a_i = 7;

    operand_b_i = 6;

    #10;

    operand_a_i = 4;

    operand_b_i = 16;

    #10;

    operand_a_i = 19;

    operand_b_i = 7;

    #10;

    operand_a_i = 4;

    operand_b_i = 5;

    #10;

    operand_a_i = 2;

    operand_b_i = 4;

    #10;

    operand_a_i = 6;

    operand_b_i = 1;

    #10;

    operand_a_i = 13;

    operand_b_i = 1;

    #10;

    operand_a_i = 2;

    operand_b_i = 7;

    #10;

    operand_a_i = 5;

    operand_b_i = 19;

    #10;

    operand_a_i = 17;

    operand_b_i = 19;

    #10;

    operand_a_i = 20;

    operand_b_i = 11;

    #10;

    operand_a_i = 12;

    operand_b_i = 15;

    #10;

    operand_a_i = 14;

    operand_b_i = 7;

    #10;

    operand_a_i = 7;

    operand_b_i = 12;

    #10;

    operand_a_i = 15;

    operand_b_i = 5;

    #10;

    operand_a_i = 11;

    operand_b_i = 6;

    #10;

    operand_a_i = 8;

    operand_b_i = 5;

    #10;

    operand_a_i = 2;

    operand_b_i = 17;

    #10;

    operand_a_i = 8;

    operand_b_i = 13;

    #10;

    operand_a_i = 5;

    operand_b_i = 3;

    #10;

    operand_a_i = 13;

    operand_b_i = 9;

    #10;

    operand_a_i = 4;

    operand_b_i = 10;

    #10;

    operand_a_i = 15;

    operand_b_i = 7;

    #10;

    operand_a_i = 18;

    operand_b_i = 17;

    #10;

    operand_a_i = 4;

    operand_b_i = 20;

    #10;

    operand_a_i = 12;

    operand_b_i = 14;

    #10;

    operand_a_i = 13;

    operand_b_i = 12;

    #10;

    operand_a_i = 15;

    operand_b_i = 14;

    #10;

    operand_a_i = 16;

    operand_b_i = 12;

    #10;

    operand_a_i = 2;

    operand_b_i = 4;

    #10;

    operand_a_i = 19;

    operand_b_i = 20;

    #10;

    operand_a_i = 15;

    operand_b_i = 17;

    #10;

    operand_a_i = 8;

    operand_b_i = 13;

    #10;

    operand_a_i = 6;

    operand_b_i = 3;

    #10;

    operand_a_i = 16;

    operand_b_i = 12;

    #10;

    operand_a_i = 1;

    operand_b_i = 4;

    #10;

    operand_a_i = 3;

    operand_b_i = 17;

    #10;

    operand_a_i = 16;

    operand_b_i = 13;

    #10;

    operand_a_i = 16;

    operand_b_i = 13;

    #10;

    operand_a_i = 13;

    operand_b_i = 2;

    #10;

    operand_a_i = 13;

    operand_b_i = 9;

    #10;

    operand_a_i = 10;

    operand_b_i = 3;

    #10;

    operand_a_i = 17;

    operand_b_i = 1;

    #10;

    operand_a_i = 19;

    operand_b_i = 12;

    #10;

    operand_a_i = 11;

    operand_b_i = 1;

    #10;

    operand_a_i = 14;

    operand_b_i = 4;

    #10;

    operand_a_i = 2;

    operand_b_i = 20;

    #10;

    operand_a_i = 8;

    operand_b_i = 11;

    #10;

    operand_a_i = 15;

    operand_b_i = 14;

    #10;

    operand_a_i = 17;

    operand_b_i = 12;

    #10;

    operand_a_i = 12;

    operand_b_i = 11;

    #10;

    operand_a_i = 2;

    operand_b_i = 13;

    #10;

    operand_a_i = 3;

    operand_b_i = 15;

    #10;

    operand_a_i = 9;

    operand_b_i = 14;

    #10;

    operand_a_i = 15;

    operand_b_i = 11;

    #10;

    operand_a_i = 11;

    operand_b_i = 20;

    #10;

    operand_a_i = 17;

    operand_b_i = 4;

    #10;

    operand_a_i = 4;

    operand_b_i = 3;

    #10;

    operand_a_i = 9;

    operand_b_i = 2;

    #10;

    operand_a_i = 17;

    operand_b_i = 9;

    #10;

    operand_a_i = 4;

    operand_b_i = 10;

    #10;

    operand_a_i = 18;

    operand_b_i = 16;

    #10;

    operand_a_i = 4;

    operand_b_i = 14;

    #10;

    operand_a_i = 8;

    operand_b_i = 19;

    #10;

    operand_a_i = 16;

    operand_b_i = 19;

    #10;

    operand_a_i = 17;

    operand_b_i = 2;

    #10;

    operand_a_i = 8;

    operand_b_i = 6;

    #10;

    operand_a_i = 3;

    operand_b_i = 14;

    #10;

    operand_a_i = 9;

    operand_b_i = 20;

    #10;

    operand_a_i = 7;

    operand_b_i = 11;

    #10;

    operand_a_i = 17;

    operand_b_i = 19;

    #10;

    operand_a_i = 10;

    operand_b_i = 18;

    #10;

    operand_a_i = 2;

    operand_b_i = 3;

    #10;

    operand_a_i = 11;

    operand_b_i = 8;

    #10;

    operand_a_i = 19;

    operand_b_i = 20;

    #10;

    operand_a_i = 14;

    operand_b_i = 17;

    #10;

    operand_a_i = 12;

    operand_b_i = 15;

    #10;

    operand_a_i = 16;

    operand_b_i = 11;

    #10;

    operand_a_i = 4;

    operand_b_i = 9;

    #10;

    operand_a_i = 6;

    operand_b_i = 18;

    #10;

    operand_a_i = 15;

    operand_b_i = 3;

    #10;

    operand_a_i = 6;

    operand_b_i = 4;

    #10;

    operand_a_i = 7;

    operand_b_i = 1;

    #10;

    operand_a_i = 18;

    operand_b_i = 19;

    #10;

    operand_a_i = 9;

    operand_b_i = 17;

    #10;

    operand_a_i = 12;

    operand_b_i = 14;

    #10;

    operand_a_i = 4;

    operand_b_i = 12;

    #10;

    operand_a_i = 7;

    operand_b_i = 5;

    #10;

    operand_a_i = 7;

    operand_b_i = 13;

    #10;

    operand_a_i = 12;

    operand_b_i = 20;

    #10;

    operand_a_i = 20;

    operand_b_i = 5;

    #10;

    operand_a_i = 9;

    operand_b_i = 19;

    #10;

    operand_a_i = 6;

    operand_b_i = 18;

    #10;

    operand_a_i = 2;

    operand_b_i = 1;

    #10;

    operand_a_i = 9;

    operand_b_i = 8;

    #10;

    operand_a_i = 7;

    operand_b_i = 20;

    #10;

    operand_a_i = 20;

    operand_b_i = 4;

    #10;

    operand_a_i = 13;

    operand_b_i = 2;

    #10;

    operand_a_i = 1;

    operand_b_i = 8;

    #10;

    operand_a_i = 10;

    operand_b_i = 12;

    #10;

    operand_a_i = 8;

    operand_b_i = 1;

    #10;

    operand_a_i = 1;

    operand_b_i = 17;

    #10;

    operand_a_i = 14;

    operand_b_i = 4;

    #10;

    operand_a_i = 20;

    operand_b_i = 4;

    #10;

    operand_a_i = 15;

    operand_b_i = 9;

    #10;

    operand_a_i = 1;

    operand_b_i = 19;

    #10;

    operand_a_i = 11;

    operand_b_i = 6;

    #10;

    operand_a_i = 10;

    operand_b_i = 4;

    #10;

    operand_a_i = 9;

    operand_b_i = 20;

    #10;

    operand_a_i = 2;

    operand_b_i = 16;

    #10;

    operand_a_i = 13;

    operand_b_i = 5;

    #10;

    operand_a_i = 15;

    operand_b_i = 4;

    #10;

    operand_a_i = 9;

    operand_b_i = 11;

    #10;

    operand_a_i = 2;

    operand_b_i = 19;

    #10;

    operand_a_i = 6;

    operand_b_i = 8;

    #10;

    operand_a_i = 14;

    operand_b_i = 16;

    #10;

    operand_a_i = 2;

    operand_b_i = 12;

    #10;

    operand_a_i = 3;

    operand_b_i = 7;

    #10;

    operand_a_i = 1;

    operand_b_i = 9;

    #10;

    operand_a_i = 14;

    operand_b_i = 9;

    #10;

    operand_a_i = 12;

    operand_b_i = 3;

    #10;

    operand_a_i = 10;

    operand_b_i = 6;

    #10;

    operand_a_i = 18;

    operand_b_i = 15;

    #10;

    operand_a_i = 14;

    operand_b_i = 6;

    #10;

    operand_a_i = 9;

    operand_b_i = 15;

    #10;

    operand_a_i = 8;

    operand_b_i = 1;

    #10;

    operand_a_i = 15;

    operand_b_i = 7;

    #10;

    operand_a_i = 18;

    operand_b_i = 6;

    #10;

    operand_a_i = 17;

    operand_b_i = 13;

    #10;

    operand_a_i = 19;

    operand_b_i = 13;

    #10;

    operand_a_i = 10;

    operand_b_i = 12;

    #10;

    operand_a_i = 13;

    operand_b_i = 16;

    #10;

    operand_a_i = 10;

    operand_b_i = 4;

    #10;

    operand_a_i = 8;

    operand_b_i = 19;

    #10;

    operand_a_i = 14;

    operand_b_i = 20;

    #10;

    operand_a_i = 11;

    operand_b_i = 7;

    #10;

    operand_a_i = 1;

    operand_b_i = 11;

    #10;

    operand_a_i = 19;

    operand_b_i = 14;

    #10;

    operand_a_i = 18;

    operand_b_i = 3;

    #10;

    operand_a_i = 7;

    operand_b_i = 18;

    #10;

    operand_a_i = 15;

    operand_b_i = 8;

    #10;

    operand_a_i = 20;

    operand_b_i = 5;

    #10;

    operand_a_i = 5;

    operand_b_i = 19;

    #10;

    operand_a_i = 6;

    operand_b_i = 15;

    #10;

    operand_a_i = 13;

    operand_b_i = 3;

    #10;

    operand_a_i = 8;

    operand_b_i = 14;

    #10;

    operand_a_i = 15;

    operand_b_i = 7;

    #10;

    operand_a_i = 13;

    operand_b_i = 19;

    #10;

    operand_a_i = 14;

    operand_b_i = 4;

    #10;

    operand_a_i = 4;

    operand_b_i = 15;

    #10;

    operand_a_i = 17;

    operand_b_i = 20;

    #10;

    operand_a_i = 9;

    operand_b_i = 11;

    #10;

    operand_a_i = 15;

    operand_b_i = 19;

    #10;

    operand_a_i = 4;

    operand_b_i = 20;

    #10;

    operand_a_i = 13;

    operand_b_i = 12;

    #10;

    operand_a_i = 19;

    operand_b_i = 7;

    #10;

    operand_a_i = 3;

    operand_b_i = 17;

    #10;

    operand_a_i = 3;

    operand_b_i = 16;

    #10;

    operand_a_i = 18;

    operand_b_i = 19;

    #10;

    operand_a_i = 18;

    operand_b_i = 4;

    #10;

    operand_a_i = 18;

    operand_b_i = 5;

    #10;

    operand_a_i = 17;

    operand_b_i = 15;

    #10;

    operand_a_i = 3;

    operand_b_i = 2;

    #10;

    operand_a_i = 17;

    operand_b_i = 10;

    #10;

    operand_a_i = 3;

    operand_b_i = 16;

    #10;

    operand_a_i = 3;

    operand_b_i = 2;

    #10;

    operand_a_i = 11;

    operand_b_i = 18;

    #10;

    operand_a_i = 16;

    operand_b_i = 17;

    #10;

    operand_a_i = 15;

    operand_b_i = 4;

    #10;

    operand_a_i = 19;

    operand_b_i = 15;

    #10;

    operand_a_i = 6;

    operand_b_i = 5;

    #10;

    operand_a_i = 18;

    operand_b_i = 14;

    #10;

    operand_a_i = 17;

    operand_b_i = 15;

    #10;

    operand_a_i = 8;

    operand_b_i = 17;

    #10;

    operand_a_i = 8;

    operand_b_i = 9;

    #10;

    operand_a_i = 12;

    operand_b_i = 9;

    #10;

    operand_a_i = 7;

    operand_b_i = 19;

    #10;

    operand_a_i = 3;

    operand_b_i = 20;

    #10;

    operand_a_i = 10;

    operand_b_i = 11;

    #10;

    operand_a_i = 11;

    operand_b_i = 20;

    #10;

    operand_a_i = 7;

    operand_b_i = 19;

    #10;

    operand_a_i = 18;

    operand_b_i = 6;

    #10;

    operand_a_i = 4;

    operand_b_i = 6;

    #10;

    operand_a_i = 12;

    operand_b_i = 15;

    #10;

    operand_a_i = 9;

    operand_b_i = 11;

    #10;

    operand_a_i = 2;

    operand_b_i = 17;

    #10;

    operand_a_i = 8;

    operand_b_i = 18;

    #10;

    operand_a_i = 7;

    operand_b_i = 11;

    #10;

    operand_a_i = 12;

    operand_b_i = 11;

    #10;

    operand_a_i = 5;

    operand_b_i = 3;

    #10;

    operand_a_i = 17;

    operand_b_i = 4;

    #10;

    operand_a_i = 6;

    operand_b_i = 9;

    #10;

    operand_a_i = 2;

    operand_b_i = 10;

    #10;

    operand_a_i = 13;

    operand_b_i = 7;

    #10;

    operand_a_i = 6;

    operand_b_i = 20;

    #10;

    operand_a_i = 20;

    operand_b_i = 12;

    #10;

    operand_a_i = 9;

    operand_b_i = 3;

    #10;

    operand_a_i = 18;

    operand_b_i = 3;

    #10;

    operand_a_i = 7;

    operand_b_i = 12;

    #10;

    operand_a_i = 14;

    operand_b_i = 18;

    #10;

    operand_a_i = 4;

    operand_b_i = 7;

    #10;

    operand_a_i = 14;

    operand_b_i = 8;

    #10;

    operand_a_i = 6;

    operand_b_i = 14;

    #10;

    operand_a_i = 17;

    operand_b_i = 19;

    #10;

    operand_a_i = 10;

    operand_b_i = 12;

    #10;

    operand_a_i = 7;

    operand_b_i = 19;

    #10;

    operand_a_i = 7;

    operand_b_i = 8;

    #10;

    operand_a_i = 3;

    operand_b_i = 10;

    #10;

    operand_a_i = 15;

    operand_b_i = 11;

    #10;

    operand_a_i = 15;

    operand_b_i = 18;

    #10;

    operand_a_i = 3;

    operand_b_i = 7;

    #10;

    operand_a_i = 4;

    operand_b_i = 14;

    #10;

    operand_a_i = 7;

    operand_b_i = 6;

    #10;

    operand_a_i = 12;

    operand_b_i = 2;

    #10;

    operand_a_i = 13;

    operand_b_i = 5;

    #10;

    operand_a_i = 13;

    operand_b_i = 14;

    #10;

    operand_a_i = 20;

    operand_b_i = 12;

    #10;

    operand_a_i = 2;

    operand_b_i = 13;

    #10;

    operand_a_i = 2;

    operand_b_i = 12;

    #10;

    operand_a_i = 9;

    operand_b_i = 18;

    #10;

    operand_a_i = 17;

    operand_b_i = 11;

    #10;

    operand_a_i = 2;

    operand_b_i = 4;

    #10;

    operand_a_i = 17;

    operand_b_i = 18;

    #10;

    operand_a_i = 4;

    operand_b_i = 6;

    #10;

    operand_a_i = 7;

    operand_b_i = 14;

    #10;

    operand_a_i = 18;

    operand_b_i = 12;

    #10;

    operand_a_i = 6;

    operand_b_i = 11;

    #10;

    operand_a_i = 5;

    operand_b_i = 6;

    #10;

    operand_a_i = 1;

    operand_b_i = 6;

    #10;

    operand_a_i = 13;

    operand_b_i = 18;

    #10;

    operand_a_i = 3;

    operand_b_i = 1;

    #10;

    operand_a_i = 15;

    operand_b_i = 14;

    #10;

    operand_a_i = 7;

    operand_b_i = 9;

    #10;

    operand_a_i = 14;

    operand_b_i = 11;

    #10;

    operand_a_i = 4;

    operand_b_i = 10;

    #10;

    operand_a_i = 10;

    operand_b_i = 3;

    #10;

    operand_a_i = 12;

    operand_b_i = 4;

    #10;

    operand_a_i = 19;

    operand_b_i = 2;

    #10;

    operand_a_i = 6;

    operand_b_i = 4;

    #10;

    operand_a_i = 16;

    operand_b_i = 19;

    #10;

    operand_a_i = 3;

    operand_b_i = 11;

    #10;

    operand_a_i = 11;

    operand_b_i = 20;

    #10;

    operand_a_i = 18;

    operand_b_i = 20;

    #10;

    operand_a_i = 12;

    operand_b_i = 16;

    #10;

    operand_a_i = 16;

    operand_b_i = 4;

    #10;

    operand_a_i = 2;

    operand_b_i = 11;

    #10;

    operand_a_i = 19;

    operand_b_i = 6;

    #10;

    operand_a_i = 1;

    operand_b_i = 11;

    #10;

    operand_a_i = 20;

    operand_b_i = 6;

    #10;

    operand_a_i = 18;

    operand_b_i = 15;

    #10;

    operand_a_i = 13;

    operand_b_i = 11;

    #10;

    operand_a_i = 15;

    operand_b_i = 7;

    #10;

    operand_a_i = 16;

    operand_b_i = 13;

    #10;

    operand_a_i = 10;

    operand_b_i = 13;

    #10;

    operand_a_i = 4;

    operand_b_i = 1;

    #10;

    operand_a_i = 7;

    operand_b_i = 9;

    #10;

    operand_a_i = 19;

    operand_b_i = 7;

    #10;

    operand_a_i = 6;

    operand_b_i = 18;

    #10;

    operand_a_i = 11;

    operand_b_i = 2;

    #10;

    operand_a_i = 6;

    operand_b_i = 5;

    #10;

    operand_a_i = 3;

    operand_b_i = 2;

    #10;

    operand_a_i = 9;

    operand_b_i = 15;

    #10;

    operand_a_i = 11;

    operand_b_i = 12;

    #10;

    operand_a_i = 5;

    operand_b_i = 4;

    #10;

    operand_a_i = 6;

    operand_b_i = 19;

    #10;

    operand_a_i = 3;

    operand_b_i = 16;

    #10;

    operand_a_i = 18;

    operand_b_i = 3;

    #10;

    operand_a_i = 2;

    operand_b_i = 4;

    #10;

    operand_a_i = 19;

    operand_b_i = 7;

    #10;

    operand_a_i = 1;

    operand_b_i = 18;

    #10;

    operand_a_i = 2;

    operand_b_i = 15;

    #10;

    operand_a_i = 16;

    operand_b_i = 8;

    #10;

    operand_a_i = 12;

    operand_b_i = 15;

    #10;

    operand_a_i = 6;

    operand_b_i = 10;

    #10;

    operand_a_i = 6;

    operand_b_i = 13;

    #10;

    operand_a_i = 10;

    operand_b_i = 6;

    #10;

    operand_a_i = 6;

    operand_b_i = 19;

    #10;

    operand_a_i = 1;

    operand_b_i = 3;

    #10;

    operand_a_i = 13;

    operand_b_i = 12;

    #10;

    operand_a_i = 18;

    operand_b_i = 17;

    #10;

    operand_a_i = 16;

    operand_b_i = 20;

    #10;

    operand_a_i = 16;

    operand_b_i = 1;

    #10;

    operand_a_i = 15;

    operand_b_i = 16;

    #10;

    operand_a_i = 16;

    operand_b_i = 4;

    #10;

    operand_a_i = 16;

    operand_b_i = 9;

    #10;

    operand_a_i = 15;

    operand_b_i = 11;

    #10;

    operand_a_i = 2;

    operand_b_i = 7;

    #10;

    operand_a_i = 11;

    operand_b_i = 8;

    #10;

    operand_a_i = 2;

    operand_b_i = 4;

    #10;

    operand_a_i = 8;

    operand_b_i = 18;

    #10;

    operand_a_i = 11;

    operand_b_i = 14;

    #10;

    operand_a_i = 3;

    operand_b_i = 8;

    #10;

    operand_a_i = 4;

    operand_b_i = 17;

    #10;

    operand_a_i = 18;

    operand_b_i = 14;

    #10;

    operand_a_i = 7;

    operand_b_i = 9;

    #10;

    operand_a_i = 2;

    operand_b_i = 19;

    #10;

    operand_a_i = 2;

    operand_b_i = 9;

    #10;

    operand_a_i = 16;

    operand_b_i = 2;

    #10;

    operand_a_i = 13;

    operand_b_i = 12;

    #10;

    operand_a_i = 12;

    operand_b_i = 18;

    #10;

    operand_a_i = 9;

    operand_b_i = 2;

    #10;

    operand_a_i = 14;

    operand_b_i = 6;

    #10;

    operand_a_i = 2;

    operand_b_i = 12;

    #10;

    operand_a_i = 7;

    operand_b_i = 19;

    #10;

    operand_a_i = 1;

    operand_b_i = 20;

    #10;

    operand_a_i = 14;

    operand_b_i = 6;

    #10;

    operand_a_i = 18;

    operand_b_i = 14;

    #10;

    operand_a_i = 20;

    operand_b_i = 8;

    #10;

    operand_a_i = 19;

    operand_b_i = 9;

    #10;

    operand_a_i = 14;

    operand_b_i = 16;

    #10;

    operand_a_i = 8;

    operand_b_i = 19;

    #10;

    operand_a_i = 11;

    operand_b_i = 18;

    #10;

    operand_a_i = 13;

    operand_b_i = 3;

    #10;

    operand_a_i = 8;

    operand_b_i = 18;

    #10;

    operand_a_i = 14;

    operand_b_i = 20;

    #10;

    operand_a_i = 17;

    operand_b_i = 16;

    #10;

    operand_a_i = 3;

    operand_b_i = 2;

    #10;

    operand_a_i = 20;

    operand_b_i = 19;

    #10;

    operand_a_i = 5;

    operand_b_i = 17;

    #10;

    operand_a_i = 6;

    operand_b_i = 5;

    #10;

    operand_a_i = 5;

    operand_b_i = 13;

    #10;

    operand_a_i = 4;

    operand_b_i = 20;

    #10;

    operand_a_i = 4;

    operand_b_i = 8;

    #10;

    operand_a_i = 17;

    operand_b_i = 6;

    #10;

    operand_a_i = 3;

    operand_b_i = 18;

    #10;

    operand_a_i = 16;

    operand_b_i = 10;

    #10;

    operand_a_i = 10;

    operand_b_i = 5;

    #10;

    operand_a_i = 14;

    operand_b_i = 19;

    #10;

    operand_a_i = 4;

    operand_b_i = 20;

    #10;

    operand_a_i = 10;

    operand_b_i = 11;

    #10;

    operand_a_i = 11;

    operand_b_i = 12;

    #10;

    operand_a_i = 8;

    operand_b_i = 12;

    #10;

    operand_a_i = 19;

    operand_b_i = 1;

    #10;

    operand_a_i = 15;

    operand_b_i = 13;

    #10;

    operand_a_i = 4;

    operand_b_i = 16;

    #10;

    operand_a_i = 16;

    operand_b_i = 9;

    #10;

    operand_a_i = 13;

    operand_b_i = 10;

    #10;

    operand_a_i = 15;

    operand_b_i = 10;

    #10;

    operand_a_i = 4;

    operand_b_i = 15;

    #10;

    operand_a_i = 4;

    operand_b_i = 8;

    #10;

    operand_a_i = 9;

    operand_b_i = 8;

    #10;

    operand_a_i = 7;

    operand_b_i = 11;

    #10;

    operand_a_i = 8;

    operand_b_i = 9;

    #10;

    operand_a_i = 6;

    operand_b_i = 13;

    #10;

    operand_a_i = 8;

    operand_b_i = 20;

    #10;

    operand_a_i = 10;

    operand_b_i = 5;

    #10;

    operand_a_i = 4;

    operand_b_i = 11;

    #10;

    operand_a_i = 3;

    operand_b_i = 19;

    #10;

    operand_a_i = 6;

    operand_b_i = 16;

    #10;

    operand_a_i = 12;

    operand_b_i = 10;

    #10;

    operand_a_i = 3;

    operand_b_i = 17;

    #10;

    operand_a_i = 9;

    operand_b_i = 4;

    #10;

    operand_a_i = 8;

    operand_b_i = 6;

    #10;

    operand_a_i = 8;

    operand_b_i = 10;

    #10;

    operand_a_i = 1;

    operand_b_i = 16;

    #10;

    operand_a_i = 18;

    operand_b_i = 16;

    #10;

    operand_a_i = 9;

    operand_b_i = 19;

    #10;

    operand_a_i = 17;

    operand_b_i = 15;

    #10;

    operand_a_i = 7;

    operand_b_i = 9;

    #10;

    operand_a_i = 17;

    operand_b_i = 16;

    #10;

    operand_a_i = 17;

    operand_b_i = 14;

    #10;

    operand_a_i = 16;

    operand_b_i = 20;

    #10;

    operand_a_i = 13;

    operand_b_i = 6;

    #10;

    operand_a_i = 1;

    operand_b_i = 3;

    #10;

    operand_a_i = 16;

    operand_b_i = 4;

    #10;

    operand_a_i = 1;

    operand_b_i = 19;

    #10;

    operand_a_i = 5;

    operand_b_i = 19;

    #10;

    operand_a_i = 17;

    operand_b_i = 15;

    #10;

    operand_a_i = 5;

    operand_b_i = 8;

    #10;

    operand_a_i = 15;

    operand_b_i = 20;

    #10;

    operand_a_i = 11;

    operand_b_i = 13;

    #10;

    operand_a_i = 17;

    operand_b_i = 14;

    #10;

    operand_a_i = 17;

    operand_b_i = 20;

    #10;

    operand_a_i = 2;

    operand_b_i = 19;

    #10;

    operand_a_i = 17;

    operand_b_i = 2;

    #10;

    operand_a_i = 6;

    operand_b_i = 20;

    #10;

    operand_a_i = 13;

    operand_b_i = 2;

    #10;

    operand_a_i = 14;

    operand_b_i = 1;

    #10;

    operand_a_i = 20;

    operand_b_i = 18;

    #10;

    operand_a_i = 12;

    operand_b_i = 16;

    #10;

    operand_a_i = 14;

    operand_b_i = 11;

    #10;

    operand_a_i = 3;

    operand_b_i = 14;

    #10;

    operand_a_i = 3;

    operand_b_i = 7;

    #10;

    operand_a_i = 1;

    operand_b_i = 20;

    #10;

    operand_a_i = 11;

    operand_b_i = 14;

    #10;

    operand_a_i = 11;

    operand_b_i = 4;

    #10;

    operand_a_i = 2;

    operand_b_i = 4;

    #10;

    operand_a_i = 16;

    operand_b_i = 13;

    #10;

    operand_a_i = 16;

    operand_b_i = 5;

    #10;

    operand_a_i = 3;

    operand_b_i = 4;

    #10;

    operand_a_i = 15;

    operand_b_i = 16;

    #10;

    operand_a_i = 18;

    operand_b_i = 14;

    #10;

    operand_a_i = 19;

    operand_b_i = 7;

    #10;

    operand_a_i = 6;

    operand_b_i = 14;

    #10;

    operand_a_i = 16;

    operand_b_i = 18;

    #10;

    operand_a_i = 11;

    operand_b_i = 14;

    #10;

    operand_a_i = 9;

    operand_b_i = 7;

    #10;

    operand_a_i = 2;

    operand_b_i = 17;

    #10;

    operand_a_i = 20;

    operand_b_i = 6;

    #10;

    operand_a_i = 20;

    operand_b_i = 7;

    #10;

    operand_a_i = 20;

    operand_b_i = 5;

    #10;

    operand_a_i = 11;

    operand_b_i = 4;

    #10;

    operand_a_i = 2;

    operand_b_i = 16;

    #10;

    operand_a_i = 6;

    operand_b_i = 5;

    #10;

    operand_a_i = 2;

    operand_b_i = 16;

    #10;

    operand_a_i = 13;

    operand_b_i = 2;

    #10;

    operand_a_i = 10;

    operand_b_i = 16;

    #10;

    operand_a_i = 18;

    operand_b_i = 16;

    #10;

    operand_a_i = 4;

    operand_b_i = 19;

    #10;

    operand_a_i = 18;

    operand_b_i = 4;

    #10;

    operand_a_i = 16;

    operand_b_i = 2;

    #10;

    operand_a_i = 6;

    operand_b_i = 4;

    #10;

    operand_a_i = 9;

    operand_b_i = 3;

    #10;

    operand_a_i = 20;

    operand_b_i = 13;

    #10;

    operand_a_i = 3;

    operand_b_i = 11;

    #10;

    operand_a_i = 5;

    operand_b_i = 2;

    #10;

    operand_a_i = 11;

    operand_b_i = 14;

    #10;

    operand_a_i = 9;

    operand_b_i = 12;

    #10;

    operand_a_i = 17;

    operand_b_i = 18;

    #10;

    operand_a_i = 12;

    operand_b_i = 4;

    #10;

    operand_a_i = 20;

    operand_b_i = 10;

    #10;

    operand_a_i = 10;

    operand_b_i = 12;

    #10;

    operand_a_i = 5;

    operand_b_i = 17;

    #10;

    operand_a_i = 1;

    operand_b_i = 20;

    #10;

    operand_a_i = 10;

    operand_b_i = 1;

    #10;

    operand_a_i = 15;

    operand_b_i = 20;

    #10;

    operand_a_i = 14;

    operand_b_i = 5;

    #10;

    operand_a_i = 20;

    operand_b_i = 12;

    #10;

    operand_a_i = 6;

    operand_b_i = 4;

    #10;

    operand_a_i = 9;

    operand_b_i = 17;

    #10;

    operand_a_i = 3;

    operand_b_i = 7;

    #10;

    operand_a_i = 1;

    operand_b_i = 9;

    #10;

    operand_a_i = 10;

    operand_b_i = 9;

    #10;

    operand_a_i = 12;

    operand_b_i = 14;

    #10;

    operand_a_i = 6;

    operand_b_i = 15;

    #10;

    operand_a_i = 10;

    operand_b_i = 15;

    #10;

    operand_a_i = 20;

    operand_b_i = 2;

    #10;

    operand_a_i = 8;

    operand_b_i = 5;

    #10;

    operand_a_i = 5;

    operand_b_i = 12;

    #10;

    operand_a_i = 6;

    operand_b_i = 13;

    #10;

    operand_a_i = 1;

    operand_b_i = 5;

    #10;

    operand_a_i = 9;

    operand_b_i = 5;

    #10;

    operand_a_i = 12;

    operand_b_i = 5;

    #10;

    operand_a_i = 10;

    operand_b_i = 16;

    #10;

    operand_a_i = 12;

    operand_b_i = 14;

    #10;

    operand_a_i = 6;

    operand_b_i = 5;

    #10;

    operand_a_i = 20;

    operand_b_i = 5;

    #10;

    operand_a_i = 19;

    operand_b_i = 8;

    #10;

    operand_a_i = 11;

    operand_b_i = 14;

    #10;

    operand_a_i = 18;

    operand_b_i = 11;

    #10;

    operand_a_i = 13;

    operand_b_i = 20;

    #10;

    operand_a_i = 2;

    operand_b_i = 16;

    #10;

    operand_a_i = 18;

    operand_b_i = 3;

    #10;

    operand_a_i = 17;

    operand_b_i = 7;

    #10;

    operand_a_i = 19;

    operand_b_i = 20;

    #10;

    operand_a_i = 6;

    operand_b_i = 14;

    #10;

    operand_a_i = 1;

    operand_b_i = 7;

    #10;

    operand_a_i = 16;

    operand_b_i = 18;

    #10;

    operand_a_i = 10;

    operand_b_i = 11;

    #10;

    operand_a_i = 3;

    operand_b_i = 12;

    #10;

    operand_a_i = 2;

    operand_b_i = 10;

    #10;

    operand_a_i = 4;

    operand_b_i = 14;

    #10;

    operand_a_i = 11;

    operand_b_i = 10;

    #10;

    operand_a_i = 4;

    operand_b_i = 11;

    #10;

    operand_a_i = 12;

    operand_b_i = 18;

    #10;

    operand_a_i = 7;

    operand_b_i = 6;

    #10;

    operand_a_i = 13;

    operand_b_i = 19;

    #10;

    operand_a_i = 16;

    operand_b_i = 1;

    #10;

    operand_a_i = 17;

    operand_b_i = 18;

    #10;

    operand_a_i = 9;

    operand_b_i = 12;

    #10;

    operand_a_i = 10;

    operand_b_i = 17;

    #10;

    operand_a_i = 14;

    operand_b_i = 6;

    #10;

    operand_a_i = 17;

    operand_b_i = 1;

    #10;

    operand_a_i = 13;

    operand_b_i = 14;

    #10;

    operand_a_i = 7;

    operand_b_i = 3;

    #10;

    operand_a_i = 18;

    operand_b_i = 5;

    #10;

    operand_a_i = 13;

    operand_b_i = 6;

    #10;

    operand_a_i = 5;

    operand_b_i = 9;

    #10;

    operand_a_i = 9;

    operand_b_i = 6;

    #10;

    operand_a_i = 20;

    operand_b_i = 11;

    #10;

    operand_a_i = 15;

    operand_b_i = 9;

    #10;

    operand_a_i = 19;

    operand_b_i = 17;

    #10;

    operand_a_i = 6;

    operand_b_i = 18;

    #10;

    operand_a_i = 5;

    operand_b_i = 10;

    #10;

    operand_a_i = 8;

    operand_b_i = 11;

    #10;

    operand_a_i = 10;

    operand_b_i = 2;

    #10;

    operand_a_i = 16;

    operand_b_i = 20;

    #10;

    operand_a_i = 17;

    operand_b_i = 14;

    #10;

    operand_a_i = 13;

    operand_b_i = 1;

    #10;

    operand_a_i = 16;

    operand_b_i = 12;

    #10;

    operand_a_i = 10;

    operand_b_i = 8;

    #10;

    operand_a_i = 19;

    operand_b_i = 11;

    #10;

    operand_a_i = 9;

    operand_b_i = 2;

    #10;

    operand_a_i = 14;

    operand_b_i = 6;

    #10;

    operand_a_i = 20;

    operand_b_i = 7;

    #10;

    operand_a_i = 16;

    operand_b_i = 14;

    #10;

    operand_a_i = 5;

    operand_b_i = 8;

    #10;

    operand_a_i = 18;

    operand_b_i = 2;

    #10;

    operand_a_i = 19;

    operand_b_i = 9;

    #10;

    operand_a_i = 10;

    operand_b_i = 16;

    #10;

    operand_a_i = 7;

    operand_b_i = 13;

    #10;

    operand_a_i = 9;

    operand_b_i = 16;

    #10;

    operand_a_i = 6;

    operand_b_i = 12;

    #10;

    operand_a_i = 13;

    operand_b_i = 7;

    #10;

    operand_a_i = 15;

    operand_b_i = 17;

    #10;

    operand_a_i = 6;

    operand_b_i = 7;

    #10;

    operand_a_i = 6;

    operand_b_i = 7;

    #10;

    operand_a_i = 8;

    operand_b_i = 1;

    #10;

    operand_a_i = 13;

    operand_b_i = 14;

    #10;

    operand_a_i = 11;

    operand_b_i = 20;

    #10;

    operand_a_i = 19;

    operand_b_i = 1;

    #10;

    operand_a_i = 9;

    operand_b_i = 14;

    #10;

    operand_a_i = 6;

    operand_b_i = 17;

    #10;

    operand_a_i = 15;

    operand_b_i = 20;

    #10;

    operand_a_i = 6;

    operand_b_i = 10;

    #10;

    operand_a_i = 9;

    operand_b_i = 13;

    #10;

    operand_a_i = 7;

    operand_b_i = 14;

    #10;

    operand_a_i = 5;

    operand_b_i = 13;

    #10;

    operand_a_i = 2;

    operand_b_i = 15;

    #10;

    operand_a_i = 19;

    operand_b_i = 4;

    #10;

    operand_a_i = 17;

    operand_b_i = 5;

    #10;

    operand_a_i = 15;

    operand_b_i = 10;

    #10;

    operand_a_i = 10;

    operand_b_i = 2;

    #10;

    operand_a_i = 14;

    operand_b_i = 20;

    #10;

    operand_a_i = 10;

    operand_b_i = 13;

    #10;

    operand_a_i = 19;

    operand_b_i = 13;

    #10;

    operand_a_i = 4;

    operand_b_i = 18;

    #10;

    operand_a_i = 3;

    operand_b_i = 14;

    #10;

    operand_a_i = 7;

    operand_b_i = 2;

    #10;

    operand_a_i = 10;

    operand_b_i = 16;

    #10;

    operand_a_i = 2;

    operand_b_i = 15;

    #10;

    operand_a_i = 6;

    operand_b_i = 12;

    #10;

    operand_a_i = 5;

    operand_b_i = 11;

    #10;

    operand_a_i = 14;

    operand_b_i = 13;

    #10;

    operand_a_i = 4;

    operand_b_i = 14;

    #10;

    operand_a_i = 17;

    operand_b_i = 6;

    #10;

    operand_a_i = 13;

    operand_b_i = 5;

    #10;

    operand_a_i = 12;

    operand_b_i = 4;

    #10;

    operand_a_i = 1;

    operand_b_i = 9;

    #10;

    operand_a_i = 12;

    operand_b_i = 5;

    #10;

    operand_a_i = 20;

    operand_b_i = 7;

    #10;

    operand_a_i = 12;

    operand_b_i = 2;

    #10;

    operand_a_i = 20;

    operand_b_i = 11;

    #10;

    operand_a_i = 2;

    operand_b_i = 16;

    #10;

    operand_a_i = 16;

    operand_b_i = 2;

    #10;

    operand_a_i = 20;

    operand_b_i = 12;

    #10;

    operand_a_i = 3;

    operand_b_i = 1;

    #10;

    operand_a_i = 15;

    operand_b_i = 3;

    #10;

    operand_a_i = 7;

    operand_b_i = 18;

    #10;

    operand_a_i = 10;

    operand_b_i = 2;

    #10;

    operand_a_i = 18;

    operand_b_i = 9;

    #10;

    operand_a_i = 13;

    operand_b_i = 2;

    #10;

    operand_a_i = 5;

    operand_b_i = 13;

    #10;

    operand_a_i = 12;

    operand_b_i = 4;

    #10;

    operand_a_i = 15;

    operand_b_i = 7;

    #10;

    operand_a_i = 5;

    operand_b_i = 12;

    #10;

    operand_a_i = 8;

    operand_b_i = 1;

    #10;

    operand_a_i = 2;

    operand_b_i = 3;

    #10;

    operand_a_i = 3;

    operand_b_i = 10;

    #10;

    operand_a_i = 12;

    operand_b_i = 18;

    #10;

    operand_a_i = 13;

    operand_b_i = 1;

    #10;

    operand_a_i = 11;

    operand_b_i = 7;

    #10;

    operand_a_i = 8;

    operand_b_i = 16;

    #10;

    operand_a_i = 2;

    operand_b_i = 15;

    #10;

    operand_a_i = 20;

    operand_b_i = 12;

    #10;

    operand_a_i = 10;

    operand_b_i = 1;

    #10;

    operand_a_i = 3;

    operand_b_i = 16;

    #10;

    operand_a_i = 11;

    operand_b_i = 10;

    #10;

    operand_a_i = 11;

    operand_b_i = 15;

    #10;

    operand_a_i = 9;

    operand_b_i = 19;

    #10;

    operand_a_i = 14;

    operand_b_i = 10;

    #10;

    operand_a_i = 11;

    operand_b_i = 16;

    #10;

    operand_a_i = 18;

    operand_b_i = 3;

    #10;

    operand_a_i = 6;

    operand_b_i = 2;

    #10;

    operand_a_i = 5;

    operand_b_i = 1;

    #10;

    operand_a_i = 19;

    operand_b_i = 8;

    #10;

    operand_a_i = 18;

    operand_b_i = 6;

    #10;

    operand_a_i = 11;

    operand_b_i = 15;

    #10;

    operand_a_i = 3;

    operand_b_i = 6;

    #10;

    operand_a_i = 5;

    operand_b_i = 14;

    #10;

    operand_a_i = 18;

    operand_b_i = 11;

    #10;

    operand_a_i = 18;

    operand_b_i = 9;

    #10;

    operand_a_i = 14;

    operand_b_i = 6;

    #10;

    operand_a_i = 16;

    operand_b_i = 2;

    #10;

    operand_a_i = 14;

    operand_b_i = 12;

    #10;

    operand_a_i = 14;

    operand_b_i = 19;

    #10;

    operand_a_i = 2;

    operand_b_i = 15;

    #10;

    operand_a_i = 17;

    operand_b_i = 15;

    #10;

    operand_a_i = 4;

    operand_b_i = 10;

    #10;

    operand_a_i = 12;

    operand_b_i = 7;

    #10;

    operand_a_i = 12;

    operand_b_i = 3;

    #10;

    operand_a_i = 15;

    operand_b_i = 11;

    #10;

    operand_a_i = 10;

    operand_b_i = 7;

    #10;

    operand_a_i = 1;

    operand_b_i = 6;

    #10;

    operand_a_i = 6;

    operand_b_i = 9;

    #10;

    operand_a_i = 12;

    operand_b_i = 16;

    #10;

    operand_a_i = 16;

    operand_b_i = 11;

    #10;

    operand_a_i = 2;

    operand_b_i = 17;

    #10;

    operand_a_i = 7;

    operand_b_i = 17;

    #10;

    operand_a_i = 17;

    operand_b_i = 6;

    #10;

    operand_a_i = 7;

    operand_b_i = 1;

    #10;

    operand_a_i = 13;

    operand_b_i = 12;

    #10;

    operand_a_i = 20;

    operand_b_i = 12;

    #10;

    operand_a_i = 10;

    operand_b_i = 1;

    #10;

    operand_a_i = 2;

    operand_b_i = 17;

    #10;

    operand_a_i = 12;

    operand_b_i = 11;

    #10;

    operand_a_i = 12;

    operand_b_i = 8;

    #10;

    operand_a_i = 19;

    operand_b_i = 17;

    #10;

    operand_a_i = 5;

    operand_b_i = 1;

    #10;

    operand_a_i = 9;

    operand_b_i = 6;

    #10;

    operand_a_i = 16;

    operand_b_i = 19;

    #10;

    operand_a_i = 12;

    operand_b_i = 17;

    #10;

    operand_a_i = 6;

    operand_b_i = 10;

    #10;

    operand_a_i = 20;

    operand_b_i = 9;

    #10;

    operand_a_i = 1;

    operand_b_i = 8;

    #10;

    operand_a_i = 11;

    operand_b_i = 8;

    #10;

    operand_a_i = 4;

    operand_b_i = 6;

    #10;

    operand_a_i = 4;

    operand_b_i = 12;

    #10;

    operand_a_i = 20;

    operand_b_i = 1;

    #10;

    operand_a_i = 10;

    operand_b_i = 2;

    #10;

    operand_a_i = 11;

    operand_b_i = 16;

    #10;

    operand_a_i = 20;

    operand_b_i = 15;

    #10;

    operand_a_i = 7;

    operand_b_i = 20;

    #10;

    operand_a_i = 3;

    operand_b_i = 10;

    #10;

    operand_a_i = 6;

    operand_b_i = 20;

    #10;

    operand_a_i = 7;

    operand_b_i = 2;

    #10;

    operand_a_i = 15;

    operand_b_i = 8;

    #10;

    operand_a_i = 9;

    operand_b_i = 15;

    #10;

    operand_a_i = 5;

    operand_b_i = 18;

    #10;

    operand_a_i = 19;

    operand_b_i = 14;

    #10;

    operand_a_i = 10;

    operand_b_i = 11;

    #10;

    operand_a_i = 6;

    operand_b_i = 13;

    #10;

    operand_a_i = 20;

    operand_b_i = 9;

    #10;

    operand_a_i = 9;

    operand_b_i = 5;

    #10;

    operand_a_i = 7;

    operand_b_i = 14;

    #10;

    operand_a_i = 18;

    operand_b_i = 2;

    #10;

    operand_a_i = 10;

    operand_b_i = 15;

    #10;

    operand_a_i = 5;

    operand_b_i = 19;

    #10;

    operand_a_i = 10;

    operand_b_i = 14;

    #10;

    operand_a_i = 16;

    operand_b_i = 7;

    #10;

    operand_a_i = 3;

    operand_b_i = 17;

    #10;

    operand_a_i = 16;

    operand_b_i = 15;

    #10;

    operand_a_i = 16;

    operand_b_i = 17;

    #10;

    operand_a_i = 10;

    operand_b_i = 19;

    #10;

    operand_a_i = 8;

    operand_b_i = 15;

    #10;

    operand_a_i = 13;

    operand_b_i = 4;

    #10;

    operand_a_i = 12;

    operand_b_i = 13;

    #10;

    operand_a_i = 10;

    operand_b_i = 7;

    #10;

    operand_a_i = 16;

    operand_b_i = 1;

    #10;

    operand_a_i = 5;

    operand_b_i = 11;

    #10;

    operand_a_i = 2;

    operand_b_i = 19;

    #10;

    operand_a_i = 10;

    operand_b_i = 6;

    #10;

    operand_a_i = 4;

    operand_b_i = 16;

    #10;

    operand_a_i = 5;

    operand_b_i = 12;

    #10;

    operand_a_i = 15;

    operand_b_i = 17;

    #10;

    operand_a_i = 7;

    operand_b_i = 15;

    #10;

    operand_a_i = 12;

    operand_b_i = 10;

    #10;

    operand_a_i = 8;

    operand_b_i = 17;

    #10;

    operand_a_i = 11;

    operand_b_i = 5;

    #10;

    operand_a_i = 17;

    operand_b_i = 1;

    #10;

    operand_a_i = 8;

    operand_b_i = 19;

    #10;

    operand_a_i = 1;

    operand_b_i = 8;

    #10;

    operand_a_i = 8;

    operand_b_i = 17;

    #10;

    operand_a_i = 10;

    operand_b_i = 19;

    #10;

    operand_a_i = 2;

    operand_b_i = 18;

    #10;

    operand_a_i = 9;

    operand_b_i = 19;

    #10;

    operand_a_i = 13;

    operand_b_i = 4;

    #10;

    operand_a_i = 12;

    operand_b_i = 20;

    #10;

    operand_a_i = 2;

    operand_b_i = 12;

    #10;

    operand_a_i = 9;

    operand_b_i = 16;

    #10;

    operand_a_i = 6;

    operand_b_i = 1;

    #10;

    operand_a_i = 18;

    operand_b_i = 10;

    #10;

    operand_a_i = 1;

    operand_b_i = 8;

    #10;

    operand_a_i = 14;

    operand_b_i = 16;

    #10;

    operand_a_i = 11;

    operand_b_i = 10;

    #10;

    operand_a_i = 11;

    operand_b_i = 18;

    #10;

    operand_a_i = 8;

    operand_b_i = 11;

    #10;

    operand_a_i = 18;

    operand_b_i = 13;

    #10;

    operand_a_i = 17;

    operand_b_i = 14;

    #10;

    operand_a_i = 2;

    operand_b_i = 8;

    #10;

    operand_a_i = 1;

    operand_b_i = 16;

    #10;

    operand_a_i = 8;

    operand_b_i = 10;

    #10;

    operand_a_i = 2;

    operand_b_i = 11;

    #10;

    operand_a_i = 12;

    operand_b_i = 16;

    #10;

    operand_a_i = 18;

    operand_b_i = 5;

    #10;

    operand_a_i = 12;

    operand_b_i = 15;

    #10;

    operand_a_i = 15;

    operand_b_i = 18;

    #10;

    operand_a_i = 12;

    operand_b_i = 2;

    #10;

    operand_a_i = 15;

    operand_b_i = 12;

    #10;

    operand_a_i = 8;

    operand_b_i = 10;

    #10;

    operand_a_i = 2;

    operand_b_i = 10;

    #10;

    operand_a_i = 8;

    operand_b_i = 11;

    #10;

    operand_a_i = 7;

    operand_b_i = 1;

    #10;

    operand_a_i = 15;

    operand_b_i = 3;

    #10;

    operand_a_i = 10;

    operand_b_i = 18;

    #10;

    operand_a_i = 16;

    operand_b_i = 8;

    #10;

    operand_a_i = 17;

    operand_b_i = 11;

    #10;

    operand_a_i = 1;

    operand_b_i = 9;

    #10;

    operand_a_i = 20;

    operand_b_i = 11;

    #10;

    operand_a_i = 7;

    operand_b_i = 12;

    #10;

    operand_a_i = 7;

    operand_b_i = 14;

    #10;

    operand_a_i = 12;

    operand_b_i = 13;

    #10;

    operand_a_i = 19;

    operand_b_i = 2;

    #10;

    operand_a_i = 12;

    operand_b_i = 10;

    #10;

    operand_a_i = 4;

    operand_b_i = 13;

    #10;

    operand_a_i = 20;

    operand_b_i = 10;

    #10;

    operand_a_i = 14;

    operand_b_i = 18;

    #10;

    operand_a_i = 11;

    operand_b_i = 10;

    #10;

    operand_a_i = 4;

    operand_b_i = 10;

    #10;

    operand_a_i = 19;

    operand_b_i = 6;

    #10;

    operand_a_i = 2;

    operand_b_i = 12;

    #10;

    operand_a_i = 6;

    operand_b_i = 14;

    #10;

    operand_a_i = 4;

    operand_b_i = 7;

    #10;

    operand_a_i = 17;

    operand_b_i = 9;

    #10;

    operand_a_i = 13;

    operand_b_i = 5;

    #10;

    operand_a_i = 17;

    operand_b_i = 18;

    #10;

    operand_a_i = 19;

    operand_b_i = 9;

    #10;

    operand_a_i = 12;

    operand_b_i = 1;

    #10;

    operand_a_i = 2;

    operand_b_i = 3;

    #10;

    operand_a_i = 8;

    operand_b_i = 7;

    #10;

    operand_a_i = 7;

    operand_b_i = 18;

    #10;

    operand_a_i = 17;

    operand_b_i = 7;

    #10;

    operand_a_i = 7;

    operand_b_i = 18;

    #10;

    operand_a_i = 9;

    operand_b_i = 1;

    #10;

    operand_a_i = 9;

    operand_b_i = 5;

    #10;

    operand_a_i = 12;

    operand_b_i = 16;

    #10;

    operand_a_i = 20;

    operand_b_i = 2;

    #10;

    operand_a_i = 12;

    operand_b_i = 16;

    #10;

    operand_a_i = 2;

    operand_b_i = 5;

    #10;

    operand_a_i = 20;

    operand_b_i = 15;

    #10;

    operand_a_i = 4;

    operand_b_i = 19;

    #10;

    operand_a_i = 3;

    operand_b_i = 17;

    #10;

    operand_a_i = 7;

    operand_b_i = 12;

    #10;

    operand_a_i = 10;

    operand_b_i = 15;

    #10;

    operand_a_i = 17;

    operand_b_i = 11;

    #10;

    operand_a_i = 2;

    operand_b_i = 17;

    #10;

    operand_a_i = 1;

    operand_b_i = 11;

    #10;

    operand_a_i = 12;

    operand_b_i = 8;

    #10;

    operand_a_i = 15;

    operand_b_i = 13;

    #10;

    operand_a_i = 6;

    operand_b_i = 15;

    #10;

    operand_a_i = 14;

    operand_b_i = 1;

    #10;

    operand_a_i = 2;

    operand_b_i = 5;

    #10;

    operand_a_i = 6;

    operand_b_i = 9;

    #10;

    operand_a_i = 6;

    operand_b_i = 3;

    #10;

    operand_a_i = 13;

    operand_b_i = 8;

    #10;

    operand_a_i = 16;

    operand_b_i = 17;

    #10;

    operand_a_i = 13;

    operand_b_i = 7;

    #10;

    operand_a_i = 7;

    operand_b_i = 14;

    #10;

    operand_a_i = 9;

    operand_b_i = 19;

    #10;

    operand_a_i = 15;

    operand_b_i = 13;

    #10;

    operand_a_i = 19;

    operand_b_i = 15;

    #10;

    operand_a_i = 18;

    operand_b_i = 4;

    #10;

    operand_a_i = 1;

    operand_b_i = 20;

    #10;

    operand_a_i = 10;

    operand_b_i = 9;

    #10;

    operand_a_i = 8;

    operand_b_i = 17;

    #10;

    operand_a_i = 9;

    operand_b_i = 8;

    #10;

    operand_a_i = 18;

    operand_b_i = 9;

    #10;

    operand_a_i = 14;

    operand_b_i = 3;

    #10;

    operand_a_i = 18;

    operand_b_i = 6;

    #10;

    operand_a_i = 18;

    operand_b_i = 11;

    #10;

    operand_a_i = 7;

    operand_b_i = 3;

    #10;

    operand_a_i = 1;

    operand_b_i = 12;

    #10;

    operand_a_i = 3;

    operand_b_i = 2;

    #10;

    operand_a_i = 6;

    operand_b_i = 3;

    #10;

    operand_a_i = 9;

    operand_b_i = 15;

    #10;

    operand_a_i = 6;

    operand_b_i = 16;

    #10;

    operand_a_i = 15;

    operand_b_i = 19;

    #10;

    operand_a_i = 17;

    operand_b_i = 2;

    #10;

    operand_a_i = 17;

    operand_b_i = 9;

    #10;

    operand_a_i = 8;

    operand_b_i = 3;

    #10;

    operand_a_i = 7;

    operand_b_i = 14;

    #10;

    operand_a_i = 5;

    operand_b_i = 19;

    #10;

    operand_a_i = 15;

    operand_b_i = 10;

    #10;

    operand_a_i = 15;

    operand_b_i = 9;

    #10;

    operand_a_i = 18;

    operand_b_i = 13;

    #10;

    operand_a_i = 5;

    operand_b_i = 11;

    #10;

    operand_a_i = 10;

    operand_b_i = 17;

    #10;

    operand_a_i = 12;

    operand_b_i = 20;

    #10;

    operand_a_i = 19;

    operand_b_i = 12;

    #10;

    operand_a_i = 14;

    operand_b_i = 13;

    #10;

    operand_a_i = 8;

    operand_b_i = 7;

    #10;

    operand_a_i = 16;

    operand_b_i = 17;

    #10;

    operand_a_i = 9;

    operand_b_i = 18;

    #10;

    operand_a_i = 19;

    operand_b_i = 4;

    #10;

    operand_a_i = 11;

    operand_b_i = 3;

    #10;

    operand_a_i = 15;

    operand_b_i = 20;

    #10;

    operand_a_i = 9;

    operand_b_i = 20;

    #10;

    operand_a_i = 6;

    operand_b_i = 5;

    #10;

    operand_a_i = 3;

    operand_b_i = 10;

    #10;

    operand_a_i = 15;

    operand_b_i = 2;

    #10;

    operand_a_i = 2;

    operand_b_i = 9;

    #10;

    operand_a_i = 12;

    operand_b_i = 18;

    #10;

    operand_a_i = 16;

    operand_b_i = 19;

    #10;

    operand_a_i = 5;

    operand_b_i = 16;

    #10;

    operand_a_i = 15;

    operand_b_i = 5;

    #10;

    operand_a_i = 16;

    operand_b_i = 10;

    #10;

    operand_a_i = 5;

    operand_b_i = 15;

    #10;

    operand_a_i = 7;

    operand_b_i = 17;

    #10;

    operand_a_i = 20;

    operand_b_i = 10;

    #10;

    operand_a_i = 18;

    operand_b_i = 20;

    #10;

    operand_a_i = 19;

    operand_b_i = 12;

    #10;

    operand_a_i = 2;

    operand_b_i = 10;

    #10;

    operand_a_i = 18;

    operand_b_i = 4;

    #10;

    operand_a_i = 11;

    operand_b_i = 4;

    #10;

    operand_a_i = 17;

    operand_b_i = 15;

    #10;

    operand_a_i = 2;

    operand_b_i = 11;

    #10;

    operand_a_i = 14;

    operand_b_i = 13;

    #10;

    operand_a_i = 15;

    operand_b_i = 20;

    #10;

    operand_a_i = 10;

    operand_b_i = 19;

    #10;

    operand_a_i = 16;

    operand_b_i = 5;

    #10;

    operand_a_i = 3;

    operand_b_i = 2;

    #10;

    operand_a_i = 2;

    operand_b_i = 3;

    #10;

    operand_a_i = 7;

    operand_b_i = 3;

    #10;

    operand_a_i = 9;

    operand_b_i = 11;

    #10;

    operand_a_i = 1;

    operand_b_i = 17;

    #10;

    operand_a_i = 15;

    operand_b_i = 18;

    #10;

    operand_a_i = 12;

    operand_b_i = 7;

    #10;

    operand_a_i = 7;

    operand_b_i = 2;

    #10;

    operand_a_i = 4;

    operand_b_i = 2;

    #10;

    operand_a_i = 13;

    operand_b_i = 12;

    #10;

    operand_a_i = 7;

    operand_b_i = 13;

    #10;

    operand_a_i = 11;

    operand_b_i = 9;

    #10;

    operand_a_i = 12;

    operand_b_i = 20;

    #10;

    operand_a_i = 12;

    operand_b_i = 8;

    #10;

    operand_a_i = 16;

    operand_b_i = 9;

    #10;

    operand_a_i = 6;

    operand_b_i = 10;

    #10;

    operand_a_i = 9;

    operand_b_i = 2;

    #10;

    operand_a_i = 1;

    operand_b_i = 11;

    #10;

    operand_a_i = 4;

    operand_b_i = 13;

    #10;

    operand_a_i = 8;

    operand_b_i = 7;

    #10;

    operand_a_i = 3;

    operand_b_i = 4;

    #10;

    operand_a_i = 16;

    operand_b_i = 5;

    #10;

    operand_a_i = 20;

    operand_b_i = 5;

    #10;

    operand_a_i = 19;

    operand_b_i = 10;

    #10;

    operand_a_i = 19;

    operand_b_i = 12;

    #10;

    operand_a_i = 12;

    operand_b_i = 18;

    #10;

    operand_a_i = 5;

    operand_b_i = 19;

    #10;

    operand_a_i = 3;

    operand_b_i = 15;

    #10;

    operand_a_i = 16;

    operand_b_i = 8;

    #10;

    operand_a_i = 8;

    operand_b_i = 2;

    #10;

    operand_a_i = 8;

    operand_b_i = 12;

    #10;

    operand_a_i = 16;

    operand_b_i = 14;

    #10;

    operand_a_i = 18;

    operand_b_i = 5;

    #10;

    operand_a_i = 17;

    operand_b_i = 4;

    #10;

    operand_a_i = 2;

    operand_b_i = 15;

    #10;

    operand_a_i = 15;

    operand_b_i = 5;

    #10;

    operand_a_i = 13;

    operand_b_i = 10;

    #10;

    operand_a_i = 6;

    operand_b_i = 8;

    #10;

    operand_a_i = 1;

    operand_b_i = 6;

    #10;

    operand_a_i = 16;

    operand_b_i = 18;

    #10;

    operand_a_i = 9;

    operand_b_i = 8;

    #10;

    operand_a_i = 6;

    operand_b_i = 16;

    #10;

    operand_a_i = 20;

    operand_b_i = 17;

    #10;

    operand_a_i = 8;

    operand_b_i = 18;

    #10;

    operand_a_i = 12;

    operand_b_i = 3;

    #10;

    operand_a_i = 14;

    operand_b_i = 16;

    #10;

    operand_a_i = 16;

    operand_b_i = 4;

    #10;

    operand_a_i = 8;

    operand_b_i = 3;

    #10;

    operand_a_i = 18;

    operand_b_i = 11;

    #10;

    operand_a_i = 2;

    operand_b_i = 7;

    #10;

    operand_a_i = 12;

    operand_b_i = 1;

    #10;

    operand_a_i = 8;

    operand_b_i = 17;

    #10;

    operand_a_i = 5;

    operand_b_i = 19;

    #10;

    operand_a_i = 4;

    operand_b_i = 8;

    #10;

    operand_a_i = 3;

    operand_b_i = 9;

    #10;

    operand_a_i = 3;

    operand_b_i = 6;

    #10;

    operand_a_i = 1;

    operand_b_i = 16;

    #10;

    operand_a_i = 19;

    operand_b_i = 5;

    #10;

    operand_a_i = 8;

    operand_b_i = 20;

    #10;

    operand_a_i = 14;

    operand_b_i = 7;

    #10;

    operand_a_i = 4;

    operand_b_i = 11;

    #10;

    operand_a_i = 13;

    operand_b_i = 19;

    #10;

    operand_a_i = 18;

    operand_b_i = 7;

    #10;

    operand_a_i = 17;

    operand_b_i = 14;

    #10;

    operand_a_i = 12;

    operand_b_i = 2;

    #10;

    operand_a_i = 3;

    operand_b_i = 12;

    #10;

    operand_a_i = 12;

    operand_b_i = 2;

    #10;

    operand_a_i = 2;

    operand_b_i = 15;

    #10;

    operand_a_i = 13;

    operand_b_i = 15;

    #10;

    operand_a_i = 10;

    operand_b_i = 19;

    #10;

    operand_a_i = 19;

    operand_b_i = 3;

    #10;

    operand_a_i = 12;

    operand_b_i = 4;

    #10;

    operand_a_i = 6;

    operand_b_i = 5;

    #10;

    operand_a_i = 11;

    operand_b_i = 12;

    #10;

    operand_a_i = 18;

    operand_b_i = 6;

    #10;

    operand_a_i = 4;

    operand_b_i = 12;

    #10;

    operand_a_i = 17;

    operand_b_i = 2;

    #10;

    operand_a_i = 5;

    operand_b_i = 8;

    #10;

    operand_a_i = 18;

    operand_b_i = 5;

    #10;

    operand_a_i = 4;

    operand_b_i = 10;

    #10;

    operand_a_i = 17;

    operand_b_i = 12;

    #10;

    operand_a_i = 9;

    operand_b_i = 13;

    #10;

    operand_a_i = 1;

    operand_b_i = 10;

    #10;

    operand_a_i = 17;

    operand_b_i = 3;

    #10;

    operand_a_i = 20;

    operand_b_i = 13;

    #10;

    operand_a_i = 16;

    operand_b_i = 8;

    #10;

    operand_a_i = 18;

    operand_b_i = 14;

    #10;

    operand_a_i = 17;

    operand_b_i = 1;

    #10;

    operand_a_i = 10;

    operand_b_i = 8;

    #10;

    operand_a_i = 8;

    operand_b_i = 1;

    #10;

    operand_a_i = 6;

    operand_b_i = 1;

    #10;

    operand_a_i = 17;

    operand_b_i = 8;

    #10;

    operand_a_i = 13;

    operand_b_i = 5;

    #10;

    operand_a_i = 13;

    operand_b_i = 6;

    #10;

    operand_a_i = 4;

    operand_b_i = 18;

    #10;

    operand_a_i = 16;

    operand_b_i = 13;

    #10;

    operand_a_i = 11;

    operand_b_i = 15;

    #10;

    operand_a_i = 1;

    operand_b_i = 19;

    #10;

    operand_a_i = 9;

    operand_b_i = 5;

    #10;

    operand_a_i = 17;

    operand_b_i = 14;

    #10;

    operand_a_i = 18;

    operand_b_i = 11;

    #10;

    operand_a_i = 1;

    operand_b_i = 13;

    #10;

    operand_a_i = 6;

    operand_b_i = 13;

    #10;

    operand_a_i = 18;

    operand_b_i = 19;

    #10;

    operand_a_i = 2;

    operand_b_i = 18;

    #10;

    operand_a_i = 9;

    operand_b_i = 11;

    #10;

    operand_a_i = 2;

    operand_b_i = 1;

    #10;

    operand_a_i = 12;

    operand_b_i = 9;

    #10;

    operand_a_i = 4;

    operand_b_i = 13;

    #10;

    operand_a_i = 13;

    operand_b_i = 11;

    #10;

    operand_a_i = 12;

    operand_b_i = 9;

    #10;

    operand_a_i = 4;

    operand_b_i = 17;

    #10;

    operand_a_i = 13;

    operand_b_i = 19;

    #10;

    operand_a_i = 10;

    operand_b_i = 9;

    #10;

    operand_a_i = 20;

    operand_b_i = 18;

    #10;

    operand_a_i = 5;

    operand_b_i = 8;

    #10;

    operand_a_i = 20;

    operand_b_i = 19;

    #10;

    operand_a_i = 18;

    operand_b_i = 7;

    #10;

    operand_a_i = 3;

    operand_b_i = 14;

    #10;

    operand_a_i = 15;

    operand_b_i = 7;

    #10;

    operand_a_i = 10;

    operand_b_i = 17;

    #10;

    operand_a_i = 20;

    operand_b_i = 14;

    #10;

    operand_a_i = 15;

    operand_b_i = 16;

    #10;

    operand_a_i = 8;

    operand_b_i = 3;

    #10;

    operand_a_i = 5;

    operand_b_i = 12;

    #10;

    operand_a_i = 4;

    operand_b_i = 10;

    #10;

    operand_a_i = 7;

    operand_b_i = 12;

    #10;

    operand_a_i = 10;

    operand_b_i = 7;

    #10;

    operand_a_i = 14;

    operand_b_i = 19;

    #10;

    operand_a_i = 3;

    operand_b_i = 2;

    #10;

    operand_a_i = 15;

    operand_b_i = 4;

    #10;

    operand_a_i = 9;

    operand_b_i = 15;

    #10;

    operand_a_i = 4;

    operand_b_i = 14;

    #10;

    operand_a_i = 18;

    operand_b_i = 8;

    #10;

    operand_a_i = 12;

    operand_b_i = 14;

    #10;

    operand_a_i = 9;

    operand_b_i = 2;

    #10;

    operand_a_i = 12;

    operand_b_i = 16;

    #10;

    operand_a_i = 9;

    operand_b_i = 14;

    #10;

    operand_a_i = 19;

    operand_b_i = 11;

    #10;

    operand_a_i = 16;

    operand_b_i = 1;

    #10;

    operand_a_i = 2;

    operand_b_i = 4;

    #10;

    operand_a_i = 13;

    operand_b_i = 14;

    #10;

    operand_a_i = 15;

    operand_b_i = 13;

    #10;

    operand_a_i = 12;

    operand_b_i = 20;

    #10;

    operand_a_i = 19;

    operand_b_i = 5;

    #10;

    operand_a_i = 19;

    operand_b_i = 3;

    #10;

    operand_a_i = 5;

    operand_b_i = 12;

    #10;

    operand_a_i = 13;

    operand_b_i = 12;

    #10;

    operand_a_i = 9;

    operand_b_i = 4;

    #10;

    operand_a_i = 9;

    operand_b_i = 11;

    #10;

    operand_a_i = 11;

    operand_b_i = 9;

    #10;

    operand_a_i = 16;

    operand_b_i = 13;

    #10;

    operand_a_i = 7;

    operand_b_i = 1;

    #10;

    operand_a_i = 19;

    operand_b_i = 8;

    #10;

    operand_a_i = 1;

    operand_b_i = 5;

    #10;

    operand_a_i = 18;

    operand_b_i = 5;

    #10;

    operand_a_i = 11;

    operand_b_i = 19;

    #10;

    operand_a_i = 15;

    operand_b_i = 4;

    #10;

    operand_a_i = 7;

    operand_b_i = 3;

    #10;

    operand_a_i = 18;

    operand_b_i = 14;

    #10;

    operand_a_i = 9;

    operand_b_i = 4;

    #10;

    operand_a_i = 4;

    operand_b_i = 19;

    #10;

    operand_a_i = 4;

    operand_b_i = 12;

    #10;

    operand_a_i = 13;

    operand_b_i = 11;

    #10;

    operand_a_i = 3;

    operand_b_i = 9;

    #10;

    operand_a_i = 15;

    operand_b_i = 1;

    #10;

    operand_a_i = 5;

    operand_b_i = 16;

    #10;

    operand_a_i = 12;

    operand_b_i = 15;

    #10;

    operand_a_i = 11;

    operand_b_i = 9;

    #10;

    operand_a_i = 1;

    operand_b_i = 18;

    #10;

    operand_a_i = 2;

    operand_b_i = 12;

    #10;

    operand_a_i = 7;

    operand_b_i = 16;

    #10;

    operand_a_i = 4;

    operand_b_i = 3;

    #10;

    operand_a_i = 16;

    operand_b_i = 19;

    #10;

    operand_a_i = 19;

    operand_b_i = 6;

    #10;

    operand_a_i = 2;

    operand_b_i = 11;

    #10;

    operand_a_i = 9;

    operand_b_i = 12;

    #10;

    operand_a_i = 14;

    operand_b_i = 12;

    #10;

    operand_a_i = 7;

    operand_b_i = 8;

    #10;

    operand_a_i = 2;

    operand_b_i = 5;

    #10;

    operand_a_i = 6;

    operand_b_i = 14;

    #10;

    operand_a_i = 3;

    operand_b_i = 11;

    #10;

    operand_a_i = 7;

    operand_b_i = 3;

    #10;

    operand_a_i = 20;

    operand_b_i = 9;

    #10;

    operand_a_i = 2;

    operand_b_i = 1;

    #10;

    operand_a_i = 7;

    operand_b_i = 20;

    #10;

    operand_a_i = 13;

    operand_b_i = 20;

    #10;

    operand_a_i = 14;

    operand_b_i = 6;

    #10;

    operand_a_i = 12;

    operand_b_i = 19;

    #10;

    operand_a_i = 1;

    operand_b_i = 2;

    #10;

    operand_a_i = 19;

    operand_b_i = 14;

    #10;

    operand_a_i = 1;

    operand_b_i = 8;

    #10;

    operand_a_i = 16;

    operand_b_i = 2;

    #10;

    operand_a_i = 5;

    operand_b_i = 10;

    #10;

    operand_a_i = 2;

    operand_b_i = 15;

    #10;

    operand_a_i = 15;

    operand_b_i = 14;

    #10;

    operand_a_i = 8;

    operand_b_i = 1;

    #10;

    operand_a_i = 13;

    operand_b_i = 17;

    #10;

    operand_a_i = 5;

    operand_b_i = 17;

    #10;

    operand_a_i = 14;

    operand_b_i = 5;

    #10;

    operand_a_i = 8;

    operand_b_i = 1;

    #10;

    operand_a_i = 20;

    operand_b_i = 17;

    #10;

    operand_a_i = 5;

    operand_b_i = 13;

    #10;

    operand_a_i = 6;

    operand_b_i = 3;

    #10;

    operand_a_i = 19;

    operand_b_i = 5;

    #10;

    operand_a_i = 10;

    operand_b_i = 16;

    #10;

    operand_a_i = 7;

    operand_b_i = 9;

    #10;

    operand_a_i = 16;

    operand_b_i = 7;

    #10;

    operand_a_i = 8;

    operand_b_i = 2;

    #10;

    operand_a_i = 7;

    operand_b_i = 16;

    #10;

    operand_a_i = 6;

    operand_b_i = 19;

    #10;

    operand_a_i = 8;

    operand_b_i = 2;

    #10;

    operand_a_i = 20;

    operand_b_i = 17;

    #10;

    operand_a_i = 3;

    operand_b_i = 6;

    #10;

    operand_a_i = 9;

    operand_b_i = 12;

    #10;

    operand_a_i = 2;

    operand_b_i = 13;

    #10;

    operand_a_i = 16;

    operand_b_i = 11;

    #10;

    operand_a_i = 13;

    operand_b_i = 17;

    #10;

    operand_a_i = 10;

    operand_b_i = 4;

    #10;

    operand_a_i = 3;

    operand_b_i = 1;

    #10;

    operand_a_i = 12;

    operand_b_i = 14;

    #10;

    operand_a_i = 15;

    operand_b_i = 18;

    #10;

    operand_a_i = 7;

    operand_b_i = 3;

    #10;

    operand_a_i = 6;

    operand_b_i = 16;

    #10;

    operand_a_i = 8;

    operand_b_i = 6;

    #10;

    operand_a_i = 6;

    operand_b_i = 7;

    #10;

    operand_a_i = 19;

    operand_b_i = 14;

    #10;

    operand_a_i = 9;

    operand_b_i = 7;

    #10;

    operand_a_i = 18;

    operand_b_i = 3;

    #10;

    operand_a_i = 16;

    operand_b_i = 1;

    #10;

    operand_a_i = 3;

    operand_b_i = 11;

    #10;

    operand_a_i = 9;

    operand_b_i = 18;

    #10;

    operand_a_i = 15;

    operand_b_i = 3;

    #10;

    operand_a_i = 20;

    operand_b_i = 18;

    #10;

    operand_a_i = 16;

    operand_b_i = 9;

    #10;

    operand_a_i = 14;

    operand_b_i = 16;

    #10;

    operand_a_i = 9;

    operand_b_i = 20;

    #10;

    operand_a_i = 19;

    operand_b_i = 4;

    #10;

    operand_a_i = 16;

    operand_b_i = 12;

    #10;

    operand_a_i = 19;

    operand_b_i = 10;

    #10;

    operand_a_i = 16;

    operand_b_i = 2;

    #10;

    operand_a_i = 17;

    operand_b_i = 20;

    #10;

    operand_a_i = 3;

    operand_b_i = 19;

    #10;

    operand_a_i = 9;

    operand_b_i = 6;

    #10;

    operand_a_i = 1;

    operand_b_i = 7;

    #10;

    operand_a_i = 9;

    operand_b_i = 13;

    #10;

    operand_a_i = 9;

    operand_b_i = 10;

    #10;

    operand_a_i = 12;

    operand_b_i = 16;

    #10;

    operand_a_i = 1;

    operand_b_i = 15;

    #10;

    operand_a_i = 12;

    operand_b_i = 6;

    #10;

    operand_a_i = 18;

    operand_b_i = 20;

    #10;

    operand_a_i = 14;

    operand_b_i = 10;

    #10;

    operand_a_i = 4;

    operand_b_i = 6;

    #10;

    operand_a_i = 2;

    operand_b_i = 7;

    #10;

    operand_a_i = 15;

    operand_b_i = 3;

    #10;

    operand_a_i = 8;

    operand_b_i = 16;

    #10;

    operand_a_i = 10;

    operand_b_i = 3;

    #10;

    operand_a_i = 2;

    operand_b_i = 11;

    #10;

    operand_a_i = 9;

    operand_b_i = 10;

    #10;

    operand_a_i = 13;

    operand_b_i = 16;

    #10;

    operand_a_i = 3;

    operand_b_i = 15;

    #10;

    operand_a_i = 4;

    operand_b_i = 11;

    #10;

    operand_a_i = 1;

    operand_b_i = 11;

    #10;

    operand_a_i = 17;

    operand_b_i = 14;

    #10;

    operand_a_i = 14;

    operand_b_i = 2;

    #10;

    operand_a_i = 17;

    operand_b_i = 1;

    #10;

    operand_a_i = 6;

    operand_b_i = 5;

    #10;

    operand_a_i = 4;

    operand_b_i = 1;

    #10;

    operand_a_i = 4;

    operand_b_i = 10;

    #10;

    operand_a_i = 4;

    operand_b_i = 7;

    #10;

    operand_a_i = 16;

    operand_b_i = 9;

    #10;

    operand_a_i = 19;

    operand_b_i = 15;

    #10;

    operand_a_i = 12;

    operand_b_i = 2;

    #10;

    operand_a_i = 4;

    operand_b_i = 1;

    #10;

    operand_a_i = 11;

    operand_b_i = 8;

    #10;

    operand_a_i = 4;

    operand_b_i = 3;

    #10;

    operand_a_i = 7;

    operand_b_i = 4;

    #10;

    operand_a_i = 11;

    operand_b_i = 6;

    #10;

    operand_a_i = 13;

    operand_b_i = 20;

    #10;

    operand_a_i = 9;

    operand_b_i = 7;

    #10;

    operand_a_i = 1;

    operand_b_i = 14;

    #10;

    operand_a_i = 10;

    operand_b_i = 12;

    #10;

    operand_a_i = 8;

    operand_b_i = 6;

    #10;

    operand_a_i = 2;

    operand_b_i = 12;

    #10;

    operand_a_i = 15;

    operand_b_i = 1;

    #10;

    operand_a_i = 20;

    operand_b_i = 2;

    #10;

    operand_a_i = 9;

    operand_b_i = 3;

    #10;

    operand_a_i = 1;

    operand_b_i = 4;

    #10;

    operand_a_i = 5;

    operand_b_i = 6;

    #10;

    operand_a_i = 10;

    operand_b_i = 13;

    #10;

    operand_a_i = 16;

    operand_b_i = 6;

    #10;

    operand_a_i = 9;

    operand_b_i = 14;

    #10;

    operand_a_i = 13;

    operand_b_i = 2;

    #10;

    operand_a_i = 9;

    operand_b_i = 13;

    #10;

    operand_a_i = 4;

    operand_b_i = 10;

    #10;

    operand_a_i = 4;

    operand_b_i = 1;

    #10;

    operand_a_i = 9;

    operand_b_i = 20;

    #10;

    operand_a_i = 16;

    operand_b_i = 3;

    #10;

    operand_a_i = 2;

    operand_b_i = 17;

    #10;

    operand_a_i = 13;

    operand_b_i = 1;

    #10;

    operand_a_i = 11;

    operand_b_i = 5;

    #10;

    operand_a_i = 13;

    operand_b_i = 4;

    #10;

    operand_a_i = 3;

    operand_b_i = 8;

    #10;

    operand_a_i = 6;

    operand_b_i = 3;

    #10;

    operand_a_i = 11;

    operand_b_i = 8;

    #10;

    operand_a_i = 7;

    operand_b_i = 11;

    #10;

    operand_a_i = 4;

    operand_b_i = 9;

    #10;

    operand_a_i = 11;

    operand_b_i = 9;

    #10;

    operand_a_i = 12;

    operand_b_i = 17;

    #10;

    operand_a_i = 10;

    operand_b_i = 8;

    #10;

    operand_a_i = 19;

    operand_b_i = 7;

    #10;

    operand_a_i = 11;

    operand_b_i = 12;

    #10;

    operand_a_i = 16;

    operand_b_i = 4;

    #10;

    operand_a_i = 12;

    operand_b_i = 11;

    #10;

    operand_a_i = 18;

    operand_b_i = 7;

    #10;

    operand_a_i = 4;

    operand_b_i = 9;

    #10;

    operand_a_i = 9;

    operand_b_i = 10;

    #10;

    operand_a_i = 16;

    operand_b_i = 19;

    #10;

    operand_a_i = 8;

    operand_b_i = 7;

    #10;

    operand_a_i = 9;

    operand_b_i = 15;

    #10;

    operand_a_i = 12;

    operand_b_i = 2;

    #10;

    operand_a_i = 19;

    operand_b_i = 15;

    #10;

    operand_a_i = 3;

    operand_b_i = 19;

    #10;

    operand_a_i = 5;

    operand_b_i = 11;

    #10;

    operand_a_i = 6;

    operand_b_i = 3;

    #10;

    operand_a_i = 12;

    operand_b_i = 17;

    #10;

    operand_a_i = 15;

    operand_b_i = 4;

    #10;

    operand_a_i = 15;

    operand_b_i = 20;

    #10;

    operand_a_i = 15;

    operand_b_i = 3;

    #10;

    operand_a_i = 4;

    operand_b_i = 3;

    #10;

    operand_a_i = 5;

    operand_b_i = 19;

    #10;

    operand_a_i = 4;

    operand_b_i = 14;

    #10;

    operand_a_i = 2;

    operand_b_i = 12;

    #10;

    operand_a_i = 14;

    operand_b_i = 2;

    #10;

    operand_a_i = 11;

    operand_b_i = 12;

    #10;

    operand_a_i = 20;

    operand_b_i = 8;

    #10;

    operand_a_i = 9;

    operand_b_i = 11;

    #10;

    operand_a_i = 5;

    operand_b_i = 6;

    #10;

    operand_a_i = 5;

    operand_b_i = 15;

    #10;

    operand_a_i = 5;

    operand_b_i = 13;

    #10;

    operand_a_i = 1;

    operand_b_i = 5;

    #10;

    operand_a_i = 11;

    operand_b_i = 16;

    #10;

    operand_a_i = 14;

    operand_b_i = 10;

    #10;

    operand_a_i = 8;

    operand_b_i = 14;

    #10;

    operand_a_i = 5;

    operand_b_i = 11;

    #10;

    operand_a_i = 10;

    operand_b_i = 20;

    #10;

    operand_a_i = 12;

    operand_b_i = 13;

    #10;

    operand_a_i = 5;

    operand_b_i = 18;

    #10;

    operand_a_i = 19;

    operand_b_i = 2;

    #10;

    operand_a_i = 20;

    operand_b_i = 18;

    #10;

    operand_a_i = 8;

    operand_b_i = 16;

    #10;

    operand_a_i = 17;

    operand_b_i = 16;

    #10;

    operand_a_i = 18;

    operand_b_i = 8;

    #10;

    operand_a_i = 12;

    operand_b_i = 11;

    #10;

    operand_a_i = 20;

    operand_b_i = 3;

    #10;

    operand_a_i = 13;

    operand_b_i = 15;

    #10;

    operand_a_i = 1;

    operand_b_i = 5;

    #10;

    operand_a_i = 16;

    operand_b_i = 12;

    #10;

    operand_a_i = 7;

    operand_b_i = 18;

    #10;

    operand_a_i = 5;

    operand_b_i = 7;

    #10;

    operand_a_i = 16;

    operand_b_i = 18;

    #10;

    operand_a_i = 4;

    operand_b_i = 17;

    #10;

    operand_a_i = 17;

    operand_b_i = 19;

    #10;

    operand_a_i = 14;

    operand_b_i = 13;

    #10;

    operand_a_i = 12;

    operand_b_i = 7;

    #10;

    operand_a_i = 12;

    operand_b_i = 11;

    #10;

    operand_a_i = 18;

    operand_b_i = 8;

    #10;

    operand_a_i = 14;

    operand_b_i = 9;

    #10;

    operand_a_i = 7;

    operand_b_i = 6;

    #10;

    operand_a_i = 10;

    operand_b_i = 7;

    #10;

    operand_a_i = 12;

    operand_b_i = 1;

    #10;

    operand_a_i = 2;

    operand_b_i = 7;

    #10;

    operand_a_i = 11;

    operand_b_i = 4;

    #10;

    operand_a_i = 7;

    operand_b_i = 3;

    #10;

    operand_a_i = 13;

    operand_b_i = 3;

    #10;

    operand_a_i = 6;

    operand_b_i = 9;

    #10;

    operand_a_i = 15;

    operand_b_i = 7;

    #10;

    operand_a_i = 7;

    operand_b_i = 6;

    #10;

    operand_a_i = 9;

    operand_b_i = 12;

    #10;

    operand_a_i = 15;

    operand_b_i = 13;

    #10;

    operand_a_i = 7;

    operand_b_i = 15;

    #10;

    operand_a_i = 12;

    operand_b_i = 20;

    #10;

    operand_a_i = 3;

    operand_b_i = 9;

    #10;

    operand_a_i = 7;

    operand_b_i = 2;

    #10;

    operand_a_i = 12;

    operand_b_i = 13;

    #10;

    operand_a_i = 13;

    operand_b_i = 1;

    #10;

    operand_a_i = 7;

    operand_b_i = 5;

    #10;

    $finish;
  end
endmodule
