`timescale 1ns/1ns

module test;

  logic clk;

  logic rst_n;

  logic start;

  logic [15:0] ain;

  logic [15:0] bin;

  logic [31:0] yout;

  logic done;


  // Device Under Test (DUT)

  verified_multi_16bit dut(
    .clk(clk),
    .rst_n(rst_n),
    .start(start),
    .ain(ain),
    .bin(bin),
    .yout(yout),
    .done(done)
  );


  always #5 clk = ~clk;


  initial begin

    $dumpfile("verified_multi_16bit.vcd");

    $dumpvars(0, test);

    clk = 0;

    rst_n = 0;

    start = 0;

    ain = 0;

    bin = 0;

    #15;

    ain = 13604;

    bin = 24193;

    rst_n = 1;

    start = 0;

    #5;

    ain = 13604;

    bin = 24193;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 54793;

    bin = 22115;

    rst_n = 1;

    start = 0;

    #5;

    ain = 54793;

    bin = 22115;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 31501;

    bin = 39309;

    rst_n = 1;

    start = 0;

    #5;

    ain = 31501;

    bin = 39309;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 33893;

    bin = 21010;

    rst_n = 1;

    start = 0;

    #5;

    ain = 33893;

    bin = 21010;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 58113;

    bin = 52493;

    rst_n = 1;

    start = 0;

    #5;

    ain = 58113;

    bin = 52493;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 61814;

    bin = 52541;

    rst_n = 1;

    start = 0;

    #5;

    ain = 61814;

    bin = 52541;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 22509;

    bin = 63372;

    rst_n = 1;

    start = 0;

    #5;

    ain = 22509;

    bin = 63372;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 59897;

    bin = 9414;

    rst_n = 1;

    start = 0;

    #5;

    ain = 59897;

    bin = 9414;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 33989;

    bin = 53930;

    rst_n = 1;

    start = 0;

    #5;

    ain = 33989;

    bin = 53930;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 63461;

    bin = 29303;

    rst_n = 1;

    start = 0;

    #5;

    ain = 63461;

    bin = 29303;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 54802;

    bin = 56207;

    rst_n = 1;

    start = 0;

    #5;

    ain = 54802;

    bin = 56207;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 27122;

    bin = 38606;

    rst_n = 1;

    start = 0;

    #5;

    ain = 27122;

    bin = 38606;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 31464;

    bin = 20165;

    rst_n = 1;

    start = 0;

    #5;

    ain = 31464;

    bin = 20165;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 18780;

    bin = 10429;

    rst_n = 1;

    start = 0;

    #5;

    ain = 18780;

    bin = 10429;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 22573;

    bin = 9829;

    rst_n = 1;

    start = 0;

    #5;

    ain = 22573;

    bin = 9829;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 25187;

    bin = 34570;

    rst_n = 1;

    start = 0;

    #5;

    ain = 25187;

    bin = 34570;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 8832;

    bin = 8480;

    rst_n = 1;

    start = 0;

    #5;

    ain = 8832;

    bin = 8480;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 17834;

    bin = 52381;

    rst_n = 1;

    start = 0;

    #5;

    ain = 17834;

    bin = 52381;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 16022;

    bin = 47123;

    rst_n = 1;

    start = 0;

    #5;

    ain = 16022;

    bin = 47123;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 14349;

    bin = 54867;

    rst_n = 1;

    start = 0;

    #5;

    ain = 14349;

    bin = 54867;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 56683;

    bin = 10965;

    rst_n = 1;

    start = 0;

    #5;

    ain = 56683;

    bin = 10965;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 18946;

    bin = 16046;

    rst_n = 1;

    start = 0;

    #5;

    ain = 18946;

    bin = 16046;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 59677;

    bin = 29391;

    rst_n = 1;

    start = 0;

    #5;

    ain = 59677;

    bin = 29391;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 18723;

    bin = 25866;

    rst_n = 1;

    start = 0;

    #5;

    ain = 18723;

    bin = 25866;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 2762;

    bin = 19516;

    rst_n = 1;

    start = 0;

    #5;

    ain = 2762;

    bin = 19516;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 48626;

    bin = 24970;

    rst_n = 1;

    start = 0;

    #5;

    ain = 48626;

    bin = 24970;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 45889;

    bin = 13528;

    rst_n = 1;

    start = 0;

    #5;

    ain = 45889;

    bin = 13528;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 62328;

    bin = 4745;

    rst_n = 1;

    start = 0;

    #5;

    ain = 62328;

    bin = 4745;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 3563;

    bin = 26038;

    rst_n = 1;

    start = 0;

    #5;

    ain = 3563;

    bin = 26038;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 63942;

    bin = 5038;

    rst_n = 1;

    start = 0;

    #5;

    ain = 63942;

    bin = 5038;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 700;

    bin = 56618;

    rst_n = 1;

    start = 0;

    #5;

    ain = 700;

    bin = 56618;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 39435;

    bin = 48753;

    rst_n = 1;

    start = 0;

    #5;

    ain = 39435;

    bin = 48753;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 16773;

    bin = 21839;

    rst_n = 1;

    start = 0;

    #5;

    ain = 16773;

    bin = 21839;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 24635;

    bin = 13114;

    rst_n = 1;

    start = 0;

    #5;

    ain = 24635;

    bin = 13114;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 12926;

    bin = 19221;

    rst_n = 1;

    start = 0;

    #5;

    ain = 12926;

    bin = 19221;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 39921;

    bin = 19417;

    rst_n = 1;

    start = 0;

    #5;

    ain = 39921;

    bin = 19417;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 1890;

    bin = 64332;

    rst_n = 1;

    start = 0;

    #5;

    ain = 1890;

    bin = 64332;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 21919;

    bin = 41359;

    rst_n = 1;

    start = 0;

    #5;

    ain = 21919;

    bin = 41359;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 43512;

    bin = 24759;

    rst_n = 1;

    start = 0;

    #5;

    ain = 43512;

    bin = 24759;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 22175;

    bin = 37980;

    rst_n = 1;

    start = 0;

    #5;

    ain = 22175;

    bin = 37980;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 49243;

    bin = 14217;

    rst_n = 1;

    start = 0;

    #5;

    ain = 49243;

    bin = 14217;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 12873;

    bin = 16080;

    rst_n = 1;

    start = 0;

    #5;

    ain = 12873;

    bin = 16080;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 49367;

    bin = 64593;

    rst_n = 1;

    start = 0;

    #5;

    ain = 49367;

    bin = 64593;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 12182;

    bin = 32524;

    rst_n = 1;

    start = 0;

    #5;

    ain = 12182;

    bin = 32524;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 52930;

    bin = 60872;

    rst_n = 1;

    start = 0;

    #5;

    ain = 52930;

    bin = 60872;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 23159;

    bin = 60733;

    rst_n = 1;

    start = 0;

    #5;

    ain = 23159;

    bin = 60733;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 56082;

    bin = 126;

    rst_n = 1;

    start = 0;

    #5;

    ain = 56082;

    bin = 126;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 33133;

    bin = 59193;

    rst_n = 1;

    start = 0;

    #5;

    ain = 33133;

    bin = 59193;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 36639;

    bin = 63187;

    rst_n = 1;

    start = 0;

    #5;

    ain = 36639;

    bin = 63187;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 12165;

    bin = 34936;

    rst_n = 1;

    start = 0;

    #5;

    ain = 12165;

    bin = 34936;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 22875;

    bin = 19273;

    rst_n = 1;

    start = 0;

    #5;

    ain = 22875;

    bin = 19273;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 44607;

    bin = 44842;

    rst_n = 1;

    start = 0;

    #5;

    ain = 44607;

    bin = 44842;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 25432;

    bin = 14470;

    rst_n = 1;

    start = 0;

    #5;

    ain = 25432;

    bin = 14470;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 3214;

    bin = 62108;

    rst_n = 1;

    start = 0;

    #5;

    ain = 3214;

    bin = 62108;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 39418;

    bin = 48166;

    rst_n = 1;

    start = 0;

    #5;

    ain = 39418;

    bin = 48166;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 6003;

    bin = 46243;

    rst_n = 1;

    start = 0;

    #5;

    ain = 6003;

    bin = 46243;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 43055;

    bin = 37555;

    rst_n = 1;

    start = 0;

    #5;

    ain = 43055;

    bin = 37555;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 22111;

    bin = 3396;

    rst_n = 1;

    start = 0;

    #5;

    ain = 22111;

    bin = 3396;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 65015;

    bin = 14027;

    rst_n = 1;

    start = 0;

    #5;

    ain = 65015;

    bin = 14027;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 6886;

    bin = 56154;

    rst_n = 1;

    start = 0;

    #5;

    ain = 6886;

    bin = 56154;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 49449;

    bin = 58093;

    rst_n = 1;

    start = 0;

    #5;

    ain = 49449;

    bin = 58093;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 27866;

    bin = 46693;

    rst_n = 1;

    start = 0;

    #5;

    ain = 27866;

    bin = 46693;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 58037;

    bin = 38111;

    rst_n = 1;

    start = 0;

    #5;

    ain = 58037;

    bin = 38111;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 6521;

    bin = 65348;

    rst_n = 1;

    start = 0;

    #5;

    ain = 6521;

    bin = 65348;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 3280;

    bin = 2858;

    rst_n = 1;

    start = 0;

    #5;

    ain = 3280;

    bin = 2858;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 44459;

    bin = 53006;

    rst_n = 1;

    start = 0;

    #5;

    ain = 44459;

    bin = 53006;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 44508;

    bin = 48282;

    rst_n = 1;

    start = 0;

    #5;

    ain = 44508;

    bin = 48282;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 29437;

    bin = 707;

    rst_n = 1;

    start = 0;

    #5;

    ain = 29437;

    bin = 707;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 60758;

    bin = 59726;

    rst_n = 1;

    start = 0;

    #5;

    ain = 60758;

    bin = 59726;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 30311;

    bin = 13322;

    rst_n = 1;

    start = 0;

    #5;

    ain = 30311;

    bin = 13322;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 47542;

    bin = 35384;

    rst_n = 1;

    start = 0;

    #5;

    ain = 47542;

    bin = 35384;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 34681;

    bin = 50360;

    rst_n = 1;

    start = 0;

    #5;

    ain = 34681;

    bin = 50360;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 49044;

    bin = 23955;

    rst_n = 1;

    start = 0;

    #5;

    ain = 49044;

    bin = 23955;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 11268;

    bin = 51801;

    rst_n = 1;

    start = 0;

    #5;

    ain = 11268;

    bin = 51801;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 27099;

    bin = 56909;

    rst_n = 1;

    start = 0;

    #5;

    ain = 27099;

    bin = 56909;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 47065;

    bin = 9837;

    rst_n = 1;

    start = 0;

    #5;

    ain = 47065;

    bin = 9837;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 57974;

    bin = 18890;

    rst_n = 1;

    start = 0;

    #5;

    ain = 57974;

    bin = 18890;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 11702;

    bin = 29077;

    rst_n = 1;

    start = 0;

    #5;

    ain = 11702;

    bin = 29077;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 6726;

    bin = 39684;

    rst_n = 1;

    start = 0;

    #5;

    ain = 6726;

    bin = 39684;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 25079;

    bin = 1897;

    rst_n = 1;

    start = 0;

    #5;

    ain = 25079;

    bin = 1897;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 47796;

    bin = 36232;

    rst_n = 1;

    start = 0;

    #5;

    ain = 47796;

    bin = 36232;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 55592;

    bin = 1069;

    rst_n = 1;

    start = 0;

    #5;

    ain = 55592;

    bin = 1069;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 12487;

    bin = 39982;

    rst_n = 1;

    start = 0;

    #5;

    ain = 12487;

    bin = 39982;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 58376;

    bin = 17692;

    rst_n = 1;

    start = 0;

    #5;

    ain = 58376;

    bin = 17692;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 42749;

    bin = 1833;

    rst_n = 1;

    start = 0;

    #5;

    ain = 42749;

    bin = 1833;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 36892;

    bin = 26502;

    rst_n = 1;

    start = 0;

    #5;

    ain = 36892;

    bin = 26502;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 2266;

    bin = 50749;

    rst_n = 1;

    start = 0;

    #5;

    ain = 2266;

    bin = 50749;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 42854;

    bin = 50288;

    rst_n = 1;

    start = 0;

    #5;

    ain = 42854;

    bin = 50288;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 1139;

    bin = 39354;

    rst_n = 1;

    start = 0;

    #5;

    ain = 1139;

    bin = 39354;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 45918;

    bin = 31226;

    rst_n = 1;

    start = 0;

    #5;

    ain = 45918;

    bin = 31226;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 1493;

    bin = 63002;

    rst_n = 1;

    start = 0;

    #5;

    ain = 1493;

    bin = 63002;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 185;

    bin = 24887;

    rst_n = 1;

    start = 0;

    #5;

    ain = 185;

    bin = 24887;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 14230;

    bin = 8640;

    rst_n = 1;

    start = 0;

    #5;

    ain = 14230;

    bin = 8640;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 40742;

    bin = 6838;

    rst_n = 1;

    start = 0;

    #5;

    ain = 40742;

    bin = 6838;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 33661;

    bin = 4060;

    rst_n = 1;

    start = 0;

    #5;

    ain = 33661;

    bin = 4060;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 22406;

    bin = 65400;

    rst_n = 1;

    start = 0;

    #5;

    ain = 22406;

    bin = 65400;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 39806;

    bin = 32987;

    rst_n = 1;

    start = 0;

    #5;

    ain = 39806;

    bin = 32987;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 46799;

    bin = 11129;

    rst_n = 1;

    start = 0;

    #5;

    ain = 46799;

    bin = 11129;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 58618;

    bin = 61025;

    rst_n = 1;

    start = 0;

    #5;

    ain = 58618;

    bin = 61025;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 2327;

    bin = 30881;

    rst_n = 1;

    start = 0;

    #5;

    ain = 2327;

    bin = 30881;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 37254;

    bin = 38480;

    rst_n = 1;

    start = 0;

    #5;

    ain = 37254;

    bin = 38480;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 23029;

    bin = 34869;

    rst_n = 1;

    start = 0;

    #5;

    ain = 23029;

    bin = 34869;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 35369;

    bin = 30145;

    rst_n = 1;

    start = 0;

    #5;

    ain = 35369;

    bin = 30145;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 29893;

    bin = 46232;

    rst_n = 1;

    start = 0;

    #5;

    ain = 29893;

    bin = 46232;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 31563;

    bin = 17011;

    rst_n = 1;

    start = 0;

    #5;

    ain = 31563;

    bin = 17011;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    ain = 59116;

    bin = 5770;

    rst_n = 1;

    start = 0;

    #5;

    ain = 59116;

    bin = 5770;

    rst_n = 1;

    start = 1;

    #200 rst_n = 0;

    #0 start = 0;

    #45;

    #50;

    $finish;
  end
endmodule
