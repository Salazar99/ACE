`timescale 1ns/1ns

module test;

  logic clk;

  logic [7:0] a;

  logic [7:0] b;

  logic cin;

  logic [7:0] sum;

  logic cout;


  // Device Under Test (DUT)

  verified_adder_8bit dut(
    .clk(clk),
    .a(a),
    .b(b),
    .cin(cin),
    .sum(sum),
    .cout(cout)
  );


  always #5 clk = ~clk;


  initial begin

    $dumpfile("verified_adder_8bit_eq_256.vcd");

    $dumpvars(0, test);

    clk = 0;

    a = 14;

    b = 241;

    cin = 1;

    #10;

    a = 104;

    b = 151;

    cin = 1;

    #10;

    a = 208;

    b = 47;

    cin = 1;

    #10;

    a = 238;

    b = 17;

    cin = 1;

    #10;

    a = 72;

    b = 183;

    cin = 1;

    #10;

    a = 184;

    b = 72;

    cin = 0;

    #10;

    a = 87;

    b = 168;

    cin = 1;

    #10;

    a = 229;

    b = 26;

    cin = 1;

    #10;

    a = 189;

    b = 66;

    cin = 1;

    #10;

    a = 217;

    b = 38;

    cin = 1;

    #10;

    a = 224;

    b = 31;

    cin = 1;

    #10;

    a = 234;

    b = 22;

    cin = 0;

    #10;

    a = 244;

    b = 11;

    cin = 1;

    #10;

    a = 102;

    b = 154;

    cin = 0;

    #10;

    a = 134;

    b = 122;

    cin = 0;

    #10;

    a = 81;

    b = 174;

    cin = 1;

    #10;

    a = 53;

    b = 203;

    cin = 0;

    #10;

    a = 215;

    b = 41;

    cin = 0;

    #10;

    a = 46;

    b = 210;

    cin = 0;

    #10;

    a = 53;

    b = 202;

    cin = 1;

    #10;

    a = 249;

    b = 6;

    cin = 1;

    #10;

    a = 228;

    b = 27;

    cin = 1;

    #10;

    a = 239;

    b = 16;

    cin = 1;

    #10;

    a = 161;

    b = 95;

    cin = 0;

    #10;

    a = 154;

    b = 101;

    cin = 1;

    #10;

    a = 7;

    b = 248;

    cin = 1;

    #10;

    a = 236;

    b = 20;

    cin = 0;

    #10;

    a = 76;

    b = 179;

    cin = 1;

    #10;

    a = 62;

    b = 194;

    cin = 0;

    #10;

    a = 90;

    b = 165;

    cin = 1;

    #10;

    a = 57;

    b = 199;

    cin = 0;

    #10;

    a = 52;

    b = 204;

    cin = 0;

    #10;

    a = 150;

    b = 105;

    cin = 1;

    #10;

    a = 210;

    b = 46;

    cin = 0;

    #10;

    a = 203;

    b = 53;

    cin = 0;

    #10;

    a = 0;

    b = 255;

    cin = 1;

    #10;

    a = 150;

    b = 105;

    cin = 1;

    #10;

    a = 195;

    b = 61;

    cin = 0;

    #10;

    a = 98;

    b = 158;

    cin = 0;

    #10;

    a = 239;

    b = 16;

    cin = 1;

    #10;

    a = 15;

    b = 240;

    cin = 1;

    #10;

    a = 119;

    b = 136;

    cin = 1;

    #10;

    a = 190;

    b = 66;

    cin = 0;

    #10;

    a = 141;

    b = 115;

    cin = 0;

    #10;

    a = 58;

    b = 197;

    cin = 1;

    #10;

    a = 43;

    b = 212;

    cin = 1;

    #10;

    a = 211;

    b = 45;

    cin = 0;

    #10;

    a = 16;

    b = 239;

    cin = 1;

    #10;

    a = 219;

    b = 36;

    cin = 1;

    #10;

    a = 87;

    b = 168;

    cin = 1;

    #10;

    a = 102;

    b = 154;

    cin = 0;

    #10;

    a = 2;

    b = 253;

    cin = 1;

    #10;

    a = 44;

    b = 212;

    cin = 0;

    #10;

    a = 126;

    b = 130;

    cin = 0;

    #10;

    a = 8;

    b = 248;

    cin = 0;

    #10;

    a = 244;

    b = 12;

    cin = 0;

    #10;

    a = 112;

    b = 143;

    cin = 1;

    #10;

    a = 132;

    b = 124;

    cin = 0;

    #10;

    a = 246;

    b = 10;

    cin = 0;

    #10;

    a = 2;

    b = 254;

    cin = 0;

    #10;

    a = 141;

    b = 115;

    cin = 0;

    #10;

    a = 45;

    b = 211;

    cin = 0;

    #10;

    a = 9;

    b = 247;

    cin = 0;

    #10;

    a = 221;

    b = 34;

    cin = 1;

    #10;

    a = 39;

    b = 216;

    cin = 1;

    #10;

    a = 94;

    b = 161;

    cin = 1;

    #10;

    a = 243;

    b = 13;

    cin = 0;

    #10;

    a = 24;

    b = 231;

    cin = 1;

    #10;

    a = 132;

    b = 123;

    cin = 1;

    #10;

    a = 70;

    b = 186;

    cin = 0;

    #10;

    a = 240;

    b = 15;

    cin = 1;

    #10;

    a = 25;

    b = 231;

    cin = 0;

    #10;

    a = 125;

    b = 130;

    cin = 1;

    #10;

    a = 146;

    b = 110;

    cin = 0;

    #10;

    a = 153;

    b = 102;

    cin = 1;

    #10;

    a = 1;

    b = 254;

    cin = 1;

    #10;

    a = 43;

    b = 213;

    cin = 0;

    #10;

    a = 194;

    b = 62;

    cin = 0;

    #10;

    a = 190;

    b = 66;

    cin = 0;

    #10;

    a = 189;

    b = 67;

    cin = 0;

    #10;

    a = 101;

    b = 154;

    cin = 1;

    #10;

    a = 129;

    b = 126;

    cin = 1;

    #10;

    a = 207;

    b = 48;

    cin = 1;

    #10;

    a = 83;

    b = 172;

    cin = 1;

    #10;

    a = 177;

    b = 78;

    cin = 1;

    #10;

    a = 173;

    b = 83;

    cin = 0;

    #10;

    a = 109;

    b = 147;

    cin = 0;

    #10;

    a = 252;

    b = 3;

    cin = 1;

    #10;

    a = 216;

    b = 39;

    cin = 1;

    #10;

    a = 222;

    b = 33;

    cin = 1;

    #10;

    a = 53;

    b = 203;

    cin = 0;

    #10;

    a = 236;

    b = 20;

    cin = 0;

    #10;

    a = 68;

    b = 188;

    cin = 0;

    #10;

    a = 118;

    b = 138;

    cin = 0;

    #10;

    a = 198;

    b = 57;

    cin = 1;

    #10;

    a = 177;

    b = 79;

    cin = 0;

    #10;

    a = 250;

    b = 5;

    cin = 1;

    #10;

    a = 111;

    b = 145;

    cin = 0;

    #10;

    a = 165;

    b = 90;

    cin = 1;

    #10;

    a = 115;

    b = 140;

    cin = 1;

    #10;

    a = 221;

    b = 35;

    cin = 0;

    #10;

    a = 132;

    b = 123;

    cin = 1;

    #10;

    a = 151;

    b = 104;

    cin = 1;

    #10;

    a = 134;

    b = 122;

    cin = 0;

    #10;

    a = 98;

    b = 158;

    cin = 0;

    #10;

    a = 103;

    b = 153;

    cin = 0;

    #10;

    a = 76;

    b = 179;

    cin = 1;

    #10;

    a = 167;

    b = 89;

    cin = 0;

    #10;

    a = 71;

    b = 185;

    cin = 0;

    #10;

    a = 100;

    b = 155;

    cin = 1;

    #10;

    a = 101;

    b = 155;

    cin = 0;

    #10;

    a = 85;

    b = 171;

    cin = 0;

    #10;

    a = 48;

    b = 207;

    cin = 1;

    #10;

    a = 12;

    b = 243;

    cin = 1;

    #10;

    a = 247;

    b = 8;

    cin = 1;

    #10;

    a = 189;

    b = 67;

    cin = 0;

    #10;

    a = 237;

    b = 19;

    cin = 0;

    #10;

    a = 170;

    b = 85;

    cin = 1;

    #10;

    a = 71;

    b = 184;

    cin = 1;

    #10;

    a = 163;

    b = 93;

    cin = 0;

    #10;

    a = 184;

    b = 72;

    cin = 0;

    #10;

    a = 175;

    b = 80;

    cin = 1;

    #10;

    a = 1;

    b = 255;

    cin = 0;

    #10;

    a = 152;

    b = 104;

    cin = 0;

    #10;

    a = 21;

    b = 234;

    cin = 1;

    #10;

    a = 100;

    b = 155;

    cin = 1;

    #10;

    a = 128;

    b = 128;

    cin = 0;

    #10;

    a = 26;

    b = 229;

    cin = 1;

    #10;

    a = 243;

    b = 12;

    cin = 1;

    #10;

    a = 169;

    b = 86;

    cin = 1;

    #10;

    a = 34;

    b = 222;

    cin = 0;

    #10;

    a = 20;

    b = 235;

    cin = 1;

    #10;

    a = 216;

    b = 39;

    cin = 1;

    #10;

    a = 24;

    b = 231;

    cin = 1;

    #10;

    a = 106;

    b = 150;

    cin = 0;

    #10;

    a = 232;

    b = 24;

    cin = 0;

    #10;

    a = 95;

    b = 160;

    cin = 1;

    #10;

    a = 89;

    b = 167;

    cin = 0;

    #10;

    a = 241;

    b = 14;

    cin = 1;

    #10;

    a = 127;

    b = 128;

    cin = 1;

    #10;

    a = 87;

    b = 169;

    cin = 0;

    #10;

    a = 217;

    b = 39;

    cin = 0;

    #10;

    a = 113;

    b = 143;

    cin = 0;

    #10;

    a = 82;

    b = 174;

    cin = 0;

    #10;

    a = 231;

    b = 24;

    cin = 1;

    #10;

    a = 159;

    b = 96;

    cin = 1;

    #10;

    a = 99;

    b = 156;

    cin = 1;

    #10;

    a = 133;

    b = 123;

    cin = 0;

    #10;

    a = 188;

    b = 68;

    cin = 0;

    #10;

    a = 22;

    b = 233;

    cin = 1;

    #10;

    a = 122;

    b = 134;

    cin = 0;

    #10;

    a = 184;

    b = 71;

    cin = 1;

    #10;

    a = 66;

    b = 190;

    cin = 0;

    #10;

    a = 208;

    b = 47;

    cin = 1;

    #10;

    a = 55;

    b = 200;

    cin = 1;

    #10;

    a = 175;

    b = 80;

    cin = 1;

    #10;

    a = 169;

    b = 87;

    cin = 0;

    #10;

    a = 242;

    b = 14;

    cin = 0;

    #10;

    a = 54;

    b = 202;

    cin = 0;

    #10;

    a = 12;

    b = 244;

    cin = 0;

    #10;

    a = 186;

    b = 70;

    cin = 0;

    #10;

    a = 192;

    b = 64;

    cin = 0;

    #10;

    a = 83;

    b = 172;

    cin = 1;

    #10;

    a = 161;

    b = 94;

    cin = 1;

    #10;

    a = 163;

    b = 93;

    cin = 0;

    #10;

    a = 36;

    b = 219;

    cin = 1;

    #10;

    a = 161;

    b = 95;

    cin = 0;

    #10;

    a = 102;

    b = 153;

    cin = 1;

    #10;

    a = 184;

    b = 72;

    cin = 0;

    #10;

    a = 77;

    b = 178;

    cin = 1;

    #10;

    a = 126;

    b = 129;

    cin = 1;

    #10;

    a = 149;

    b = 107;

    cin = 0;

    #10;

    a = 17;

    b = 239;

    cin = 0;

    #10;

    a = 68;

    b = 188;

    cin = 0;

    #10;

    a = 162;

    b = 93;

    cin = 1;

    #10;

    a = 77;

    b = 179;

    cin = 0;

    #10;

    a = 74;

    b = 181;

    cin = 1;

    #10;

    a = 11;

    b = 245;

    cin = 0;

    #10;

    a = 87;

    b = 168;

    cin = 1;

    #10;

    a = 146;

    b = 110;

    cin = 0;

    #10;

    a = 242;

    b = 14;

    cin = 0;

    #10;

    a = 125;

    b = 131;

    cin = 0;

    #10;

    a = 113;

    b = 142;

    cin = 1;

    #10;

    a = 101;

    b = 155;

    cin = 0;

    #10;

    a = 2;

    b = 254;

    cin = 0;

    #10;

    a = 61;

    b = 194;

    cin = 1;

    #10;

    a = 3;

    b = 253;

    cin = 0;

    #10;

    a = 239;

    b = 16;

    cin = 1;

    #10;

    a = 164;

    b = 92;

    cin = 0;

    #10;

    a = 150;

    b = 105;

    cin = 1;

    #10;

    a = 93;

    b = 163;

    cin = 0;

    #10;

    a = 112;

    b = 143;

    cin = 1;

    #10;

    a = 28;

    b = 227;

    cin = 1;

    #10;

    a = 251;

    b = 5;

    cin = 0;

    #10;

    a = 206;

    b = 49;

    cin = 1;

    #10;

    a = 202;

    b = 54;

    cin = 0;

    #10;

    a = 249;

    b = 7;

    cin = 0;

    #10;

    a = 96;

    b = 160;

    cin = 0;

    #10;

    a = 171;

    b = 84;

    cin = 1;

    #10;

    a = 148;

    b = 108;

    cin = 0;

    #10;

    a = 71;

    b = 184;

    cin = 1;

    #10;

    a = 180;

    b = 76;

    cin = 0;

    #10;

    a = 230;

    b = 26;

    cin = 0;

    #10;

    a = 195;

    b = 61;

    cin = 0;

    #10;

    a = 134;

    b = 121;

    cin = 1;

    #10;

    a = 64;

    b = 191;

    cin = 1;

    #10;

    a = 98;

    b = 158;

    cin = 0;

    #10;

    a = 174;

    b = 81;

    cin = 1;

    #10;

    a = 15;

    b = 241;

    cin = 0;

    #10;

    a = 116;

    b = 139;

    cin = 1;

    #10;

    a = 95;

    b = 160;

    cin = 1;

    #10;

    a = 133;

    b = 123;

    cin = 0;

    #10;

    a = 19;

    b = 237;

    cin = 0;

    #10;

    a = 195;

    b = 61;

    cin = 0;

    #10;

    a = 238;

    b = 17;

    cin = 1;

    #10;

    a = 220;

    b = 35;

    cin = 1;

    #10;

    a = 225;

    b = 30;

    cin = 1;

    #10;

    a = 233;

    b = 22;

    cin = 1;

    #10;

    a = 68;

    b = 187;

    cin = 1;

    #10;

    a = 242;

    b = 13;

    cin = 1;

    #10;

    a = 177;

    b = 79;

    cin = 0;

    #10;

    a = 182;

    b = 73;

    cin = 1;

    #10;

    a = 108;

    b = 148;

    cin = 0;

    #10;

    a = 245;

    b = 10;

    cin = 1;

    #10;

    a = 223;

    b = 32;

    cin = 1;

    #10;

    a = 120;

    b = 136;

    cin = 0;

    #10;

    a = 226;

    b = 29;

    cin = 1;

    #10;

    a = 51;

    b = 204;

    cin = 1;

    #10;

    a = 120;

    b = 136;

    cin = 0;

    #10;

    a = 244;

    b = 12;

    cin = 0;

    #10;

    a = 34;

    b = 221;

    cin = 1;

    #10;

    a = 159;

    b = 96;

    cin = 1;

    #10;

    a = 18;

    b = 237;

    cin = 1;

    #10;

    a = 137;

    b = 118;

    cin = 1;

    #10;

    a = 67;

    b = 188;

    cin = 1;

    #10;

    a = 1;

    b = 255;

    cin = 0;

    #10;

    a = 237;

    b = 19;

    cin = 0;

    #10;

    a = 140;

    b = 115;

    cin = 1;

    #10;

    a = 47;

    b = 208;

    cin = 1;

    #10;

    a = 78;

    b = 178;

    cin = 0;

    #10;

    a = 218;

    b = 37;

    cin = 1;

    #10;

    a = 46;

    b = 209;

    cin = 1;

    #10;

    a = 101;

    b = 155;

    cin = 0;

    #10;

    a = 5;

    b = 250;

    cin = 1;

    #10;

    a = 181;

    b = 74;

    cin = 1;

    #10;

    a = 215;

    b = 41;

    cin = 0;

    #10;

    a = 218;

    b = 37;

    cin = 1;

    #10;

    a = 83;

    b = 173;

    cin = 0;

    #10;

    a = 135;

    b = 121;

    cin = 0;

    #10;

    a = 78;

    b = 178;

    cin = 0;

    #10;

    a = 132;

    b = 124;

    cin = 0;

    #10;

    a = 46;

    b = 209;

    cin = 1;

    #10;

    a = 120;

    b = 136;

    cin = 0;

    #10;

    a = 113;

    b = 142;

    cin = 1;

    #10;

    a = 233;

    b = 23;

    cin = 0;

    #10;

    a = 244;

    b = 12;

    cin = 0;

    #10;

    a = 168;

    b = 87;

    cin = 1;

    #10;

    a = 35;

    b = 221;

    cin = 0;

    #10;

    a = 53;

    b = 202;

    cin = 1;

    #10;

    a = 2;

    b = 253;

    cin = 1;

    #10;

    a = 46;

    b = 210;

    cin = 0;

    #10;

    a = 146;

    b = 109;

    cin = 1;

    #10;

    a = 8;

    b = 247;

    cin = 1;

    #10;

    a = 224;

    b = 31;

    cin = 1;

    #10;

    a = 132;

    b = 124;

    cin = 0;

    #10;

    a = 97;

    b = 159;

    cin = 0;

    #10;

    a = 107;

    b = 149;

    cin = 0;

    #10;

    a = 84;

    b = 171;

    cin = 1;

    #10;

    a = 64;

    b = 191;

    cin = 1;

    #10;

    a = 42;

    b = 214;

    cin = 0;

    #10;

    a = 163;

    b = 92;

    cin = 1;

    #10;

    a = 153;

    b = 103;

    cin = 0;

    #10;

    a = 206;

    b = 49;

    cin = 1;

    #10;

    a = 111;

    b = 145;

    cin = 0;

    #10;

    a = 244;

    b = 11;

    cin = 1;

    #10;

    a = 108;

    b = 148;

    cin = 0;

    #10;

    a = 222;

    b = 34;

    cin = 0;

    #10;

    a = 137;

    b = 118;

    cin = 1;

    #10;

    a = 107;

    b = 148;

    cin = 1;

    #10;

    a = 206;

    b = 50;

    cin = 0;

    #10;

    a = 82;

    b = 173;

    cin = 1;

    #10;

    a = 111;

    b = 145;

    cin = 0;

    #10;

    a = 132;

    b = 124;

    cin = 0;

    #10;

    a = 249;

    b = 7;

    cin = 0;

    #10;

    a = 145;

    b = 110;

    cin = 1;

    #10;

    a = 193;

    b = 62;

    cin = 1;

    #10;

    a = 111;

    b = 144;

    cin = 1;

    #10;

    a = 12;

    b = 243;

    cin = 1;

    #10;

    a = 218;

    b = 37;

    cin = 1;

    #10;

    a = 77;

    b = 178;

    cin = 1;

    #10;

    a = 26;

    b = 230;

    cin = 0;

    #10;

    a = 190;

    b = 66;

    cin = 0;

    #10;

    a = 165;

    b = 90;

    cin = 1;

    #10;

    a = 122;

    b = 134;

    cin = 0;

    #10;

    a = 119;

    b = 137;

    cin = 0;

    #10;

    a = 101;

    b = 155;

    cin = 0;

    #10;

    a = 108;

    b = 148;

    cin = 0;

    #10;

    a = 253;

    b = 2;

    cin = 1;

    #10;

    a = 81;

    b = 174;

    cin = 1;

    #10;

    a = 9;

    b = 246;

    cin = 1;

    #10;

    a = 15;

    b = 241;

    cin = 0;

    #10;

    a = 75;

    b = 180;

    cin = 1;

    #10;

    a = 11;

    b = 245;

    cin = 0;

    #10;

    a = 240;

    b = 16;

    cin = 0;

    #10;

    a = 179;

    b = 77;

    cin = 0;

    #10;

    a = 183;

    b = 73;

    cin = 0;

    #10;

    a = 130;

    b = 126;

    cin = 0;

    #10;

    a = 161;

    b = 95;

    cin = 0;

    #10;

    a = 157;

    b = 98;

    cin = 1;

    #10;

    a = 93;

    b = 163;

    cin = 0;

    #10;

    a = 1;

    b = 255;

    cin = 0;

    #10;

    a = 218;

    b = 37;

    cin = 1;

    #10;

    a = 207;

    b = 48;

    cin = 1;

    #10;

    a = 165;

    b = 91;

    cin = 0;

    #10;

    a = 97;

    b = 159;

    cin = 0;

    #10;

    a = 28;

    b = 227;

    cin = 1;

    #10;

    a = 214;

    b = 42;

    cin = 0;

    #10;

    a = 166;

    b = 90;

    cin = 0;

    #10;

    a = 214;

    b = 42;

    cin = 0;

    #10;

    a = 157;

    b = 99;

    cin = 0;

    #10;

    a = 171;

    b = 85;

    cin = 0;

    #10;

    a = 42;

    b = 214;

    cin = 0;

    #10;

    a = 194;

    b = 61;

    cin = 1;

    #10;

    a = 197;

    b = 58;

    cin = 1;

    #10;

    a = 215;

    b = 40;

    cin = 1;

    #10;

    a = 45;

    b = 211;

    cin = 0;

    #10;

    a = 113;

    b = 143;

    cin = 0;

    #10;

    a = 56;

    b = 199;

    cin = 1;

    #10;

    a = 61;

    b = 194;

    cin = 1;

    #10;

    a = 178;

    b = 78;

    cin = 0;

    #10;

    a = 246;

    b = 10;

    cin = 0;

    #10;

    a = 148;

    b = 107;

    cin = 1;

    #10;

    a = 226;

    b = 29;

    cin = 1;

    #10;

    a = 96;

    b = 160;

    cin = 0;

    #10;

    a = 213;

    b = 43;

    cin = 0;

    #10;

    a = 134;

    b = 121;

    cin = 1;

    #10;

    a = 34;

    b = 221;

    cin = 1;

    #10;

    a = 164;

    b = 92;

    cin = 0;

    #10;

    a = 228;

    b = 27;

    cin = 1;

    #10;

    a = 233;

    b = 22;

    cin = 1;

    #10;

    a = 189;

    b = 67;

    cin = 0;

    #10;

    a = 121;

    b = 134;

    cin = 1;

    #10;

    a = 71;

    b = 184;

    cin = 1;

    #10;

    a = 46;

    b = 210;

    cin = 0;

    #10;

    a = 200;

    b = 55;

    cin = 1;

    #10;

    a = 193;

    b = 62;

    cin = 1;

    #10;

    a = 114;

    b = 142;

    cin = 0;

    #10;

    a = 226;

    b = 29;

    cin = 1;

    #10;

    a = 41;

    b = 215;

    cin = 0;

    #10;

    a = 195;

    b = 60;

    cin = 1;

    #10;

    a = 117;

    b = 139;

    cin = 0;

    #10;

    a = 102;

    b = 154;

    cin = 0;

    #10;

    a = 188;

    b = 68;

    cin = 0;

    #10;

    a = 180;

    b = 76;

    cin = 0;

    #10;

    a = 148;

    b = 108;

    cin = 0;

    #10;

    a = 53;

    b = 202;

    cin = 1;

    #10;

    a = 94;

    b = 161;

    cin = 1;

    #10;

    a = 13;

    b = 242;

    cin = 1;

    #10;

    a = 78;

    b = 178;

    cin = 0;

    #10;

    a = 99;

    b = 156;

    cin = 1;

    #10;

    a = 70;

    b = 186;

    cin = 0;

    #10;

    a = 230;

    b = 25;

    cin = 1;

    #10;

    a = 232;

    b = 23;

    cin = 1;

    #10;

    a = 16;

    b = 239;

    cin = 1;

    #10;

    a = 144;

    b = 111;

    cin = 1;

    #10;

    a = 4;

    b = 252;

    cin = 0;

    #10;

    a = 150;

    b = 105;

    cin = 1;

    #10;

    a = 202;

    b = 54;

    cin = 0;

    #10;

    a = 80;

    b = 175;

    cin = 1;

    #10;

    a = 102;

    b = 154;

    cin = 0;

    #10;

    a = 99;

    b = 157;

    cin = 0;

    #10;

    a = 27;

    b = 228;

    cin = 1;

    #10;

    a = 177;

    b = 79;

    cin = 0;

    #10;

    a = 155;

    b = 100;

    cin = 1;

    #10;

    a = 170;

    b = 86;

    cin = 0;

    #10;

    a = 133;

    b = 122;

    cin = 1;

    #10;

    a = 121;

    b = 134;

    cin = 1;

    #10;

    a = 228;

    b = 28;

    cin = 0;

    #10;

    a = 178;

    b = 78;

    cin = 0;

    #10;

    a = 155;

    b = 100;

    cin = 1;

    #10;

    a = 254;

    b = 2;

    cin = 0;

    #10;

    a = 172;

    b = 83;

    cin = 1;

    #10;

    a = 247;

    b = 8;

    cin = 1;

    #10;

    a = 102;

    b = 154;

    cin = 0;

    #10;

    a = 206;

    b = 50;

    cin = 0;

    #10;

    a = 56;

    b = 199;

    cin = 1;

    #10;

    a = 44;

    b = 211;

    cin = 1;

    #10;

    a = 30;

    b = 225;

    cin = 1;

    #10;

    a = 113;

    b = 143;

    cin = 0;

    #10;

    a = 83;

    b = 173;

    cin = 0;

    #10;

    a = 152;

    b = 104;

    cin = 0;

    #10;

    a = 4;

    b = 252;

    cin = 0;

    #10;

    a = 35;

    b = 221;

    cin = 0;

    #10;

    a = 164;

    b = 92;

    cin = 0;

    #10;

    a = 169;

    b = 86;

    cin = 1;

    #10;

    a = 131;

    b = 124;

    cin = 1;

    #10;

    a = 90;

    b = 165;

    cin = 1;

    #10;

    a = 90;

    b = 166;

    cin = 0;

    #10;

    a = 90;

    b = 165;

    cin = 1;

    #10;

    a = 36;

    b = 220;

    cin = 0;

    #10;

    a = 68;

    b = 187;

    cin = 1;

    #10;

    a = 99;

    b = 156;

    cin = 1;

    #10;

    a = 120;

    b = 136;

    cin = 0;

    #10;

    a = 14;

    b = 242;

    cin = 0;

    #10;

    a = 133;

    b = 122;

    cin = 1;

    #10;

    a = 31;

    b = 224;

    cin = 1;

    #10;

    a = 134;

    b = 121;

    cin = 1;

    #10;

    a = 16;

    b = 240;

    cin = 0;

    #10;

    a = 28;

    b = 228;

    cin = 0;

    #10;

    a = 67;

    b = 189;

    cin = 0;

    #10;

    a = 82;

    b = 174;

    cin = 0;

    #10;

    a = 109;

    b = 147;

    cin = 0;

    #10;

    a = 194;

    b = 61;

    cin = 1;

    #10;

    a = 204;

    b = 52;

    cin = 0;

    #10;

    a = 14;

    b = 241;

    cin = 1;

    #10;

    a = 201;

    b = 55;

    cin = 0;

    #10;

    a = 66;

    b = 189;

    cin = 1;

    #10;

    a = 62;

    b = 194;

    cin = 0;

    #10;

    a = 84;

    b = 172;

    cin = 0;

    #10;

    a = 176;

    b = 80;

    cin = 0;

    #10;

    a = 45;

    b = 211;

    cin = 0;

    #10;

    a = 213;

    b = 42;

    cin = 1;

    #10;

    a = 12;

    b = 243;

    cin = 1;

    #10;

    a = 81;

    b = 175;

    cin = 0;

    #10;

    a = 197;

    b = 58;

    cin = 1;

    #10;

    a = 156;

    b = 100;

    cin = 0;

    #10;

    a = 171;

    b = 85;

    cin = 0;

    #10;

    a = 157;

    b = 99;

    cin = 0;

    #10;

    a = 26;

    b = 229;

    cin = 1;

    #10;

    a = 156;

    b = 99;

    cin = 1;

    #10;

    a = 231;

    b = 24;

    cin = 1;

    #10;

    a = 40;

    b = 215;

    cin = 1;

    #10;

    a = 207;

    b = 48;

    cin = 1;

    #10;

    a = 31;

    b = 225;

    cin = 0;

    #10;

    a = 205;

    b = 51;

    cin = 0;

    #10;

    a = 241;

    b = 15;

    cin = 0;

    #10;

    a = 112;

    b = 144;

    cin = 0;

    #10;

    a = 179;

    b = 76;

    cin = 1;

    #10;

    a = 102;

    b = 153;

    cin = 1;

    #10;

    a = 38;

    b = 218;

    cin = 0;

    #10;

    a = 164;

    b = 91;

    cin = 1;

    #10;

    a = 90;

    b = 166;

    cin = 0;

    #10;

    a = 151;

    b = 104;

    cin = 1;

    #10;

    a = 129;

    b = 127;

    cin = 0;

    #10;

    a = 79;

    b = 177;

    cin = 0;

    #10;

    a = 81;

    b = 174;

    cin = 1;

    #10;

    a = 138;

    b = 118;

    cin = 0;

    #10;

    a = 115;

    b = 141;

    cin = 0;

    #10;

    a = 110;

    b = 146;

    cin = 0;

    #10;

    a = 168;

    b = 88;

    cin = 0;

    #10;

    a = 206;

    b = 49;

    cin = 1;

    #10;

    a = 185;

    b = 70;

    cin = 1;

    #10;

    a = 158;

    b = 98;

    cin = 0;

    #10;

    a = 204;

    b = 51;

    cin = 1;

    #10;

    a = 116;

    b = 140;

    cin = 0;

    #10;

    a = 27;

    b = 229;

    cin = 0;

    #10;

    a = 168;

    b = 88;

    cin = 0;

    #10;

    a = 90;

    b = 165;

    cin = 1;

    #10;

    a = 18;

    b = 238;

    cin = 0;

    #10;

    a = 111;

    b = 144;

    cin = 1;

    #10;

    a = 53;

    b = 202;

    cin = 1;

    #10;

    a = 192;

    b = 64;

    cin = 0;

    #10;

    a = 50;

    b = 205;

    cin = 1;

    #10;

    a = 228;

    b = 27;

    cin = 1;

    #10;

    a = 207;

    b = 48;

    cin = 1;

    #10;

    a = 37;

    b = 218;

    cin = 1;

    #10;

    a = 73;

    b = 183;

    cin = 0;

    #10;

    a = 67;

    b = 188;

    cin = 1;

    #10;

    a = 202;

    b = 53;

    cin = 1;

    #10;

    a = 151;

    b = 105;

    cin = 0;

    #10;

    a = 167;

    b = 88;

    cin = 1;

    #10;

    a = 176;

    b = 80;

    cin = 0;

    #10;

    a = 142;

    b = 113;

    cin = 1;

    #10;

    a = 12;

    b = 243;

    cin = 1;

    #10;

    a = 167;

    b = 89;

    cin = 0;

    #10;

    a = 165;

    b = 91;

    cin = 0;

    #10;

    a = 153;

    b = 103;

    cin = 0;

    #10;

    a = 162;

    b = 93;

    cin = 1;

    #10;

    a = 72;

    b = 183;

    cin = 1;

    #10;

    a = 158;

    b = 97;

    cin = 1;

    #10;

    a = 201;

    b = 54;

    cin = 1;

    #10;

    a = 213;

    b = 43;

    cin = 0;

    #10;

    a = 10;

    b = 245;

    cin = 1;

    #10;

    a = 69;

    b = 187;

    cin = 0;

    #10;

    a = 222;

    b = 33;

    cin = 1;

    #10;

    a = 4;

    b = 251;

    cin = 1;

    #10;

    a = 35;

    b = 221;

    cin = 0;

    #10;

    a = 67;

    b = 188;

    cin = 1;

    #10;

    a = 47;

    b = 208;

    cin = 1;

    #10;

    a = 26;

    b = 230;

    cin = 0;

    #10;

    a = 223;

    b = 33;

    cin = 0;

    #10;

    a = 16;

    b = 239;

    cin = 1;

    #10;

    a = 100;

    b = 155;

    cin = 1;

    #10;

    a = 156;

    b = 99;

    cin = 1;

    #10;

    a = 124;

    b = 132;

    cin = 0;

    #10;

    a = 43;

    b = 213;

    cin = 0;

    #10;

    a = 20;

    b = 235;

    cin = 1;

    #10;

    a = 207;

    b = 48;

    cin = 1;

    #10;

    a = 250;

    b = 6;

    cin = 0;

    #10;

    a = 251;

    b = 5;

    cin = 0;

    #10;

    a = 227;

    b = 29;

    cin = 0;

    #10;

    a = 178;

    b = 78;

    cin = 0;

    #10;

    a = 137;

    b = 119;

    cin = 0;

    #10;

    a = 227;

    b = 29;

    cin = 0;

    #10;

    a = 196;

    b = 59;

    cin = 1;

    #10;

    a = 144;

    b = 112;

    cin = 0;

    #10;

    a = 83;

    b = 173;

    cin = 0;

    #10;

    a = 98;

    b = 157;

    cin = 1;

    #10;

    a = 28;

    b = 228;

    cin = 0;

    #10;

    a = 143;

    b = 112;

    cin = 1;

    #10;

    a = 187;

    b = 68;

    cin = 1;

    #10;

    a = 148;

    b = 107;

    cin = 1;

    #10;

    a = 198;

    b = 58;

    cin = 0;

    #10;

    a = 4;

    b = 251;

    cin = 1;

    #10;

    a = 176;

    b = 80;

    cin = 0;

    #10;

    a = 89;

    b = 166;

    cin = 1;

    #10;

    a = 220;

    b = 35;

    cin = 1;

    #10;

    a = 21;

    b = 234;

    cin = 1;

    #10;

    a = 138;

    b = 118;

    cin = 0;

    #10;

    a = 51;

    b = 204;

    cin = 1;

    #10;

    a = 104;

    b = 151;

    cin = 1;

    #10;

    a = 43;

    b = 213;

    cin = 0;

    #10;

    a = 99;

    b = 157;

    cin = 0;

    #10;

    a = 173;

    b = 82;

    cin = 1;

    #10;

    a = 171;

    b = 85;

    cin = 0;

    #10;

    a = 112;

    b = 144;

    cin = 0;

    #10;

    a = 246;

    b = 10;

    cin = 0;

    #10;

    a = 203;

    b = 52;

    cin = 1;

    #10;

    a = 186;

    b = 69;

    cin = 1;

    #10;

    a = 127;

    b = 129;

    cin = 0;

    #10;

    a = 211;

    b = 45;

    cin = 0;

    #10;

    a = 250;

    b = 6;

    cin = 0;

    #10;

    a = 249;

    b = 6;

    cin = 1;

    #10;

    a = 218;

    b = 37;

    cin = 1;

    #10;

    a = 157;

    b = 98;

    cin = 1;

    #10;

    a = 169;

    b = 87;

    cin = 0;

    #10;

    a = 117;

    b = 139;

    cin = 0;

    #10;

    a = 77;

    b = 179;

    cin = 0;

    #10;

    a = 201;

    b = 55;

    cin = 0;

    #10;

    a = 77;

    b = 178;

    cin = 1;

    #10;

    a = 19;

    b = 236;

    cin = 1;

    #10;

    a = 48;

    b = 208;

    cin = 0;

    #10;

    a = 236;

    b = 20;

    cin = 0;

    #10;

    a = 210;

    b = 46;

    cin = 0;

    #10;

    a = 49;

    b = 206;

    cin = 1;

    #10;

    a = 44;

    b = 212;

    cin = 0;

    #10;

    a = 55;

    b = 201;

    cin = 0;

    #10;

    a = 94;

    b = 161;

    cin = 1;

    #10;

    a = 103;

    b = 152;

    cin = 1;

    #10;

    a = 12;

    b = 243;

    cin = 1;

    #10;

    a = 19;

    b = 236;

    cin = 1;

    #10;

    a = 148;

    b = 108;

    cin = 0;

    #10;

    a = 221;

    b = 34;

    cin = 1;

    #10;

    a = 104;

    b = 151;

    cin = 1;

    #10;

    a = 98;

    b = 158;

    cin = 0;

    #10;

    a = 141;

    b = 115;

    cin = 0;

    #10;

    a = 128;

    b = 128;

    cin = 0;

    #10;

    a = 182;

    b = 74;

    cin = 0;

    #10;

    a = 88;

    b = 168;

    cin = 0;

    #10;

    a = 118;

    b = 137;

    cin = 1;

    #10;

    a = 191;

    b = 64;

    cin = 1;

    #10;

    a = 177;

    b = 78;

    cin = 1;

    #10;

    a = 111;

    b = 144;

    cin = 1;

    #10;

    a = 32;

    b = 224;

    cin = 0;

    #10;

    a = 122;

    b = 133;

    cin = 1;

    #10;

    a = 121;

    b = 134;

    cin = 1;

    #10;

    a = 222;

    b = 34;

    cin = 0;

    #10;

    a = 100;

    b = 156;

    cin = 0;

    #10;

    a = 121;

    b = 134;

    cin = 1;

    #10;

    a = 248;

    b = 8;

    cin = 0;

    #10;

    a = 3;

    b = 253;

    cin = 0;

    #10;

    a = 29;

    b = 226;

    cin = 1;

    #10;

    a = 131;

    b = 125;

    cin = 0;

    #10;

    a = 195;

    b = 60;

    cin = 1;

    #10;

    a = 5;

    b = 250;

    cin = 1;

    #10;

    a = 187;

    b = 69;

    cin = 0;

    #10;

    a = 186;

    b = 70;

    cin = 0;

    #10;

    a = 172;

    b = 84;

    cin = 0;

    #10;

    a = 217;

    b = 38;

    cin = 1;

    #10;

    a = 50;

    b = 206;

    cin = 0;

    #10;

    a = 191;

    b = 64;

    cin = 1;

    #10;

    a = 8;

    b = 248;

    cin = 0;

    #10;

    a = 230;

    b = 26;

    cin = 0;

    #10;

    a = 191;

    b = 65;

    cin = 0;

    #10;

    a = 205;

    b = 51;

    cin = 0;

    #10;

    a = 149;

    b = 106;

    cin = 1;

    #10;

    a = 220;

    b = 36;

    cin = 0;

    #10;

    a = 120;

    b = 135;

    cin = 1;

    #10;

    a = 69;

    b = 187;

    cin = 0;

    #10;

    a = 95;

    b = 161;

    cin = 0;

    #10;

    a = 101;

    b = 155;

    cin = 0;

    #10;

    a = 142;

    b = 114;

    cin = 0;

    #10;

    a = 139;

    b = 117;

    cin = 0;

    #10;

    a = 41;

    b = 214;

    cin = 1;

    #10;

    a = 239;

    b = 16;

    cin = 1;

    #10;

    a = 87;

    b = 168;

    cin = 1;

    #10;

    a = 27;

    b = 228;

    cin = 1;

    #10;

    a = 80;

    b = 175;

    cin = 1;

    #10;

    a = 75;

    b = 180;

    cin = 1;

    #10;

    a = 197;

    b = 59;

    cin = 0;

    #10;

    a = 147;

    b = 108;

    cin = 1;

    #10;

    a = 127;

    b = 128;

    cin = 1;

    #10;

    a = 50;

    b = 205;

    cin = 1;

    #10;

    a = 130;

    b = 126;

    cin = 0;

    #10;

    a = 94;

    b = 162;

    cin = 0;

    #10;

    a = 150;

    b = 105;

    cin = 1;

    #10;

    a = 113;

    b = 143;

    cin = 0;

    #10;

    a = 44;

    b = 211;

    cin = 1;

    #10;

    a = 202;

    b = 54;

    cin = 0;

    #10;

    a = 189;

    b = 66;

    cin = 1;

    #10;

    a = 223;

    b = 33;

    cin = 0;

    #10;

    a = 7;

    b = 249;

    cin = 0;

    #10;

    a = 192;

    b = 63;

    cin = 1;

    #10;

    a = 45;

    b = 211;

    cin = 0;

    #10;

    a = 13;

    b = 242;

    cin = 1;

    #10;

    a = 231;

    b = 24;

    cin = 1;

    #10;

    a = 166;

    b = 90;

    cin = 0;

    #10;

    a = 241;

    b = 14;

    cin = 1;

    #10;

    a = 28;

    b = 227;

    cin = 1;

    #10;

    a = 95;

    b = 161;

    cin = 0;

    #10;

    a = 88;

    b = 168;

    cin = 0;

    #10;

    a = 137;

    b = 119;

    cin = 0;

    #10;

    a = 220;

    b = 35;

    cin = 1;

    #10;

    a = 176;

    b = 80;

    cin = 0;

    #10;

    a = 205;

    b = 51;

    cin = 0;

    #10;

    a = 64;

    b = 192;

    cin = 0;

    #10;

    a = 234;

    b = 22;

    cin = 0;

    #10;

    a = 201;

    b = 54;

    cin = 1;

    #10;

    a = 117;

    b = 138;

    cin = 1;

    #10;

    a = 89;

    b = 166;

    cin = 1;

    #10;

    a = 42;

    b = 214;

    cin = 0;

    #10;

    a = 1;

    b = 255;

    cin = 0;

    #10;

    a = 127;

    b = 129;

    cin = 0;

    #10;

    a = 137;

    b = 118;

    cin = 1;

    #10;

    a = 44;

    b = 212;

    cin = 0;

    #10;

    a = 5;

    b = 251;

    cin = 0;

    #10;

    a = 94;

    b = 161;

    cin = 1;

    #10;

    a = 195;

    b = 60;

    cin = 1;

    #10;

    a = 197;

    b = 58;

    cin = 1;

    #10;

    a = 86;

    b = 169;

    cin = 1;

    #10;

    a = 84;

    b = 171;

    cin = 1;

    #10;

    a = 183;

    b = 72;

    cin = 1;

    #10;

    a = 218;

    b = 37;

    cin = 1;

    #10;

    a = 22;

    b = 234;

    cin = 0;

    #10;

    a = 42;

    b = 214;

    cin = 0;

    #10;

    a = 202;

    b = 54;

    cin = 0;

    #10;

    a = 19;

    b = 236;

    cin = 1;

    #10;

    a = 226;

    b = 29;

    cin = 1;

    #10;

    a = 245;

    b = 10;

    cin = 1;

    #10;

    a = 124;

    b = 131;

    cin = 1;

    #10;

    a = 176;

    b = 80;

    cin = 0;

    #10;

    a = 91;

    b = 165;

    cin = 0;

    #10;

    a = 160;

    b = 95;

    cin = 1;

    #10;

    a = 210;

    b = 45;

    cin = 1;

    #10;

    a = 179;

    b = 77;

    cin = 0;

    #10;

    a = 240;

    b = 16;

    cin = 0;

    #10;

    a = 94;

    b = 161;

    cin = 1;

    #10;

    a = 190;

    b = 65;

    cin = 1;

    #10;

    a = 184;

    b = 71;

    cin = 1;

    #10;

    a = 197;

    b = 58;

    cin = 1;

    #10;

    a = 103;

    b = 152;

    cin = 1;

    #10;

    a = 185;

    b = 71;

    cin = 0;

    #10;

    a = 79;

    b = 176;

    cin = 1;

    #10;

    a = 48;

    b = 208;

    cin = 0;

    #10;

    a = 95;

    b = 160;

    cin = 1;

    #10;

    a = 214;

    b = 41;

    cin = 1;

    #10;

    a = 109;

    b = 147;

    cin = 0;

    #10;

    a = 247;

    b = 9;

    cin = 0;

    #10;

    a = 152;

    b = 104;

    cin = 0;

    #10;

    a = 73;

    b = 183;

    cin = 0;

    #10;

    a = 209;

    b = 47;

    cin = 0;

    #10;

    a = 238;

    b = 18;

    cin = 0;

    #10;

    a = 110;

    b = 145;

    cin = 1;

    #10;

    a = 95;

    b = 160;

    cin = 1;

    #10;

    a = 90;

    b = 166;

    cin = 0;

    #10;

    a = 252;

    b = 3;

    cin = 1;

    #10;

    a = 80;

    b = 175;

    cin = 1;

    #10;

    a = 182;

    b = 74;

    cin = 0;

    #10;

    a = 218;

    b = 37;

    cin = 1;

    #10;

    a = 4;

    b = 251;

    cin = 1;

    #10;

    a = 152;

    b = 103;

    cin = 1;

    #10;

    a = 67;

    b = 189;

    cin = 0;

    #10;

    a = 139;

    b = 117;

    cin = 0;

    #10;

    a = 79;

    b = 176;

    cin = 1;

    #10;

    a = 32;

    b = 223;

    cin = 1;

    #10;

    a = 168;

    b = 87;

    cin = 1;

    #10;

    a = 36;

    b = 220;

    cin = 0;

    #10;

    a = 58;

    b = 198;

    cin = 0;

    #10;

    a = 144;

    b = 111;

    cin = 1;

    #10;

    a = 38;

    b = 218;

    cin = 0;

    #10;

    a = 225;

    b = 30;

    cin = 1;

    #10;

    a = 2;

    b = 254;

    cin = 0;

    #10;

    a = 41;

    b = 214;

    cin = 1;

    #10;

    a = 141;

    b = 115;

    cin = 0;

    #10;

    a = 118;

    b = 138;

    cin = 0;

    #10;

    a = 162;

    b = 94;

    cin = 0;

    #10;

    a = 204;

    b = 51;

    cin = 1;

    #10;

    a = 218;

    b = 37;

    cin = 1;

    #10;

    a = 246;

    b = 9;

    cin = 1;

    #10;

    a = 213;

    b = 42;

    cin = 1;

    #10;

    a = 182;

    b = 74;

    cin = 0;

    #10;

    a = 39;

    b = 216;

    cin = 1;

    #10;

    a = 79;

    b = 177;

    cin = 0;

    #10;

    a = 214;

    b = 41;

    cin = 1;

    #10;

    a = 199;

    b = 56;

    cin = 1;

    #10;

    a = 254;

    b = 2;

    cin = 0;

    #10;

    a = 125;

    b = 130;

    cin = 1;

    #10;

    a = 252;

    b = 4;

    cin = 0;

    #10;

    a = 112;

    b = 144;

    cin = 0;

    #10;

    a = 230;

    b = 26;

    cin = 0;

    #10;

    a = 193;

    b = 62;

    cin = 1;

    #10;

    a = 11;

    b = 245;

    cin = 0;

    #10;

    a = 54;

    b = 201;

    cin = 1;

    #10;

    a = 163;

    b = 93;

    cin = 0;

    #10;

    a = 247;

    b = 8;

    cin = 1;

    #10;

    a = 32;

    b = 223;

    cin = 1;

    #10;

    a = 222;

    b = 33;

    cin = 1;

    #10;

    a = 141;

    b = 114;

    cin = 1;

    #10;

    a = 60;

    b = 196;

    cin = 0;

    #10;

    a = 46;

    b = 210;

    cin = 0;

    #10;

    a = 109;

    b = 146;

    cin = 1;

    #10;

    a = 140;

    b = 115;

    cin = 1;

    #10;

    a = 13;

    b = 242;

    cin = 1;

    #10;

    a = 193;

    b = 63;

    cin = 0;

    #10;

    a = 68;

    b = 188;

    cin = 0;

    #10;

    a = 160;

    b = 95;

    cin = 1;

    #10;

    a = 247;

    b = 8;

    cin = 1;

    #10;

    a = 234;

    b = 22;

    cin = 0;

    #10;

    a = 55;

    b = 200;

    cin = 1;

    #10;

    a = 241;

    b = 15;

    cin = 0;

    #10;

    a = 65;

    b = 190;

    cin = 1;

    #10;

    a = 47;

    b = 209;

    cin = 0;

    #10;

    a = 114;

    b = 142;

    cin = 0;

    #10;

    a = 68;

    b = 187;

    cin = 1;

    #10;

    a = 128;

    b = 128;

    cin = 0;

    #10;

    a = 60;

    b = 196;

    cin = 0;

    #10;

    a = 64;

    b = 191;

    cin = 1;

    #10;

    a = 246;

    b = 10;

    cin = 0;

    #10;

    a = 98;

    b = 158;

    cin = 0;

    #10;

    a = 227;

    b = 28;

    cin = 1;

    #10;

    a = 136;

    b = 119;

    cin = 1;

    #10;

    a = 7;

    b = 249;

    cin = 0;

    #10;

    a = 78;

    b = 177;

    cin = 1;

    #10;

    a = 113;

    b = 142;

    cin = 1;

    #10;

    a = 87;

    b = 168;

    cin = 1;

    #10;

    a = 210;

    b = 46;

    cin = 0;

    #10;

    a = 68;

    b = 187;

    cin = 1;

    #10;

    a = 4;

    b = 252;

    cin = 0;

    #10;

    a = 118;

    b = 137;

    cin = 1;

    #10;

    a = 133;

    b = 123;

    cin = 0;

    #10;

    a = 193;

    b = 62;

    cin = 1;

    #10;

    a = 250;

    b = 6;

    cin = 0;

    #10;

    a = 69;

    b = 187;

    cin = 0;

    #10;

    a = 157;

    b = 98;

    cin = 1;

    #10;

    a = 216;

    b = 40;

    cin = 0;

    #10;

    a = 167;

    b = 89;

    cin = 0;

    #10;

    a = 217;

    b = 38;

    cin = 1;

    #10;

    a = 164;

    b = 91;

    cin = 1;

    #10;

    a = 102;

    b = 153;

    cin = 1;

    #10;

    a = 202;

    b = 54;

    cin = 0;

    #10;

    a = 53;

    b = 202;

    cin = 1;

    #10;

    a = 86;

    b = 170;

    cin = 0;

    #10;

    a = 51;

    b = 204;

    cin = 1;

    #10;

    a = 171;

    b = 84;

    cin = 1;

    #10;

    a = 93;

    b = 163;

    cin = 0;

    #10;

    a = 133;

    b = 122;

    cin = 1;

    #10;

    a = 223;

    b = 32;

    cin = 1;

    #10;

    a = 105;

    b = 151;

    cin = 0;

    #10;

    a = 42;

    b = 213;

    cin = 1;

    #10;

    a = 63;

    b = 192;

    cin = 1;

    #10;

    a = 72;

    b = 184;

    cin = 0;

    #10;

    a = 49;

    b = 207;

    cin = 0;

    #10;

    a = 233;

    b = 22;

    cin = 1;

    #10;

    a = 238;

    b = 18;

    cin = 0;

    #10;

    a = 179;

    b = 76;

    cin = 1;

    #10;

    a = 224;

    b = 31;

    cin = 1;

    #10;

    a = 84;

    b = 172;

    cin = 0;

    #10;

    a = 115;

    b = 140;

    cin = 1;

    #10;

    a = 215;

    b = 41;

    cin = 0;

    #10;

    a = 148;

    b = 107;

    cin = 1;

    #10;

    a = 35;

    b = 220;

    cin = 1;

    #10;

    a = 182;

    b = 74;

    cin = 0;

    #10;

    a = 193;

    b = 63;

    cin = 0;

    #10;

    a = 119;

    b = 137;

    cin = 0;

    #10;

    a = 145;

    b = 110;

    cin = 1;

    #10;

    a = 12;

    b = 243;

    cin = 1;

    #10;

    a = 63;

    b = 192;

    cin = 1;

    #10;

    a = 43;

    b = 213;

    cin = 0;

    #10;

    a = 39;

    b = 217;

    cin = 0;

    #10;

    a = 143;

    b = 112;

    cin = 1;

    #10;

    a = 204;

    b = 51;

    cin = 1;

    #10;

    a = 112;

    b = 143;

    cin = 1;

    #10;

    a = 155;

    b = 100;

    cin = 1;

    #10;

    a = 131;

    b = 125;

    cin = 0;

    #10;

    a = 221;

    b = 34;

    cin = 1;

    #10;

    a = 33;

    b = 223;

    cin = 0;

    #10;

    a = 226;

    b = 29;

    cin = 1;

    #10;

    a = 103;

    b = 153;

    cin = 0;

    #10;

    a = 222;

    b = 33;

    cin = 1;

    #10;

    a = 120;

    b = 136;

    cin = 0;

    #10;

    a = 93;

    b = 163;

    cin = 0;

    #10;

    a = 193;

    b = 62;

    cin = 1;

    #10;

    a = 195;

    b = 60;

    cin = 1;

    #10;

    a = 11;

    b = 244;

    cin = 1;

    #10;

    a = 34;

    b = 221;

    cin = 1;

    #10;

    a = 19;

    b = 236;

    cin = 1;

    #10;

    a = 253;

    b = 2;

    cin = 1;

    #10;

    a = 64;

    b = 191;

    cin = 1;

    #10;

    a = 89;

    b = 166;

    cin = 1;

    #10;

    a = 142;

    b = 113;

    cin = 1;

    #10;

    a = 119;

    b = 136;

    cin = 1;

    #10;

    a = 155;

    b = 100;

    cin = 1;

    #10;

    a = 81;

    b = 175;

    cin = 0;

    #10;

    a = 238;

    b = 17;

    cin = 1;

    #10;

    a = 131;

    b = 125;

    cin = 0;

    #10;

    a = 195;

    b = 60;

    cin = 1;

    #10;

    a = 164;

    b = 91;

    cin = 1;

    #10;

    a = 48;

    b = 208;

    cin = 0;

    #10;

    a = 5;

    b = 250;

    cin = 1;

    #10;

    a = 122;

    b = 134;

    cin = 0;

    #10;

    a = 77;

    b = 179;

    cin = 0;

    #10;

    a = 191;

    b = 64;

    cin = 1;

    #10;

    a = 110;

    b = 145;

    cin = 1;

    #10;

    a = 187;

    b = 69;

    cin = 0;

    #10;

    a = 19;

    b = 236;

    cin = 1;

    #10;

    a = 196;

    b = 59;

    cin = 1;

    #10;

    a = 219;

    b = 36;

    cin = 1;

    #10;

    a = 18;

    b = 237;

    cin = 1;

    #10;

    a = 170;

    b = 85;

    cin = 1;

    #10;

    a = 234;

    b = 21;

    cin = 1;

    #10;

    a = 221;

    b = 34;

    cin = 1;

    #10;

    a = 175;

    b = 81;

    cin = 0;

    #10;

    a = 172;

    b = 84;

    cin = 0;

    #10;

    a = 202;

    b = 53;

    cin = 1;

    #10;

    a = 240;

    b = 15;

    cin = 1;

    #10;

    a = 218;

    b = 37;

    cin = 1;

    #10;

    a = 97;

    b = 159;

    cin = 0;

    #10;

    a = 252;

    b = 4;

    cin = 0;

    #10;

    a = 73;

    b = 183;

    cin = 0;

    #10;

    a = 77;

    b = 178;

    cin = 1;

    #10;

    a = 30;

    b = 226;

    cin = 0;

    #10;

    a = 216;

    b = 40;

    cin = 0;

    #10;

    a = 67;

    b = 189;

    cin = 0;

    #10;

    a = 107;

    b = 149;

    cin = 0;

    #10;

    a = 233;

    b = 23;

    cin = 0;

    #10;

    a = 158;

    b = 98;

    cin = 0;

    #10;

    a = 233;

    b = 23;

    cin = 0;

    #10;

    a = 219;

    b = 37;

    cin = 0;

    #10;

    a = 50;

    b = 205;

    cin = 1;

    #10;

    a = 193;

    b = 62;

    cin = 1;

    #10;

    a = 5;

    b = 250;

    cin = 1;

    #10;

    a = 136;

    b = 120;

    cin = 0;

    #10;

    a = 38;

    b = 217;

    cin = 1;

    #10;

    a = 204;

    b = 51;

    cin = 1;

    #10;

    a = 1;

    b = 255;

    cin = 0;

    #10;

    a = 223;

    b = 32;

    cin = 1;

    #10;

    a = 144;

    b = 112;

    cin = 0;

    #10;

    a = 131;

    b = 124;

    cin = 1;

    #10;

    a = 227;

    b = 28;

    cin = 1;

    #10;

    a = 198;

    b = 57;

    cin = 1;

    #10;

    a = 43;

    b = 213;

    cin = 0;

    #10;

    a = 130;

    b = 125;

    cin = 1;

    #10;

    a = 174;

    b = 81;

    cin = 1;

    #10;

    a = 81;

    b = 174;

    cin = 1;

    #10;

    a = 83;

    b = 172;

    cin = 1;

    #10;

    a = 39;

    b = 216;

    cin = 1;

    #10;

    a = 210;

    b = 46;

    cin = 0;

    #10;

    a = 248;

    b = 7;

    cin = 1;

    #10;

    a = 209;

    b = 47;

    cin = 0;

    #10;

    a = 108;

    b = 148;

    cin = 0;

    #10;

    a = 82;

    b = 174;

    cin = 0;

    #10;

    a = 190;

    b = 65;

    cin = 1;

    #10;

    a = 46;

    b = 210;

    cin = 0;

    #10;

    a = 54;

    b = 201;

    cin = 1;

    #10;

    a = 174;

    b = 82;

    cin = 0;

    #10;

    a = 14;

    b = 242;

    cin = 0;

    #10;

    a = 239;

    b = 17;

    cin = 0;

    #10;

    a = 38;

    b = 218;

    cin = 0;

    #10;

    a = 2;

    b = 254;

    cin = 0;

    #10;

    a = 165;

    b = 91;

    cin = 0;

    #10;

    a = 40;

    b = 215;

    cin = 1;

    #10;

    a = 251;

    b = 5;

    cin = 0;

    #10;

    a = 120;

    b = 135;

    cin = 1;

    #10;

    a = 11;

    b = 245;

    cin = 0;

    #10;

    a = 77;

    b = 179;

    cin = 0;

    #10;

    a = 221;

    b = 35;

    cin = 0;

    #10;

    a = 59;

    b = 196;

    cin = 1;

    #10;

    a = 156;

    b = 100;

    cin = 0;

    #10;

    a = 114;

    b = 141;

    cin = 1;

    #10;

    a = 94;

    b = 161;

    cin = 1;

    #10;

    a = 225;

    b = 31;

    cin = 0;

    #10;

    a = 222;

    b = 34;

    cin = 0;

    #10;

    a = 169;

    b = 87;

    cin = 0;

    #10;

    a = 189;

    b = 66;

    cin = 1;

    #10;

    a = 70;

    b = 185;

    cin = 1;

    #10;

    a = 155;

    b = 100;

    cin = 1;

    #10;

    a = 34;

    b = 221;

    cin = 1;

    #10;

    a = 116;

    b = 140;

    cin = 0;

    #10;

    a = 68;

    b = 188;

    cin = 0;

    #10;

    a = 217;

    b = 39;

    cin = 0;

    #10;

    a = 172;

    b = 83;

    cin = 1;

    #10;

    a = 71;

    b = 185;

    cin = 0;

    #10;

    a = 1;

    b = 254;

    cin = 1;

    #10;

    a = 41;

    b = 214;

    cin = 1;

    #10;

    a = 170;

    b = 86;

    cin = 0;

    #10;

    a = 42;

    b = 213;

    cin = 1;

    #10;

    a = 229;

    b = 27;

    cin = 0;

    #10;

    a = 71;

    b = 184;

    cin = 1;

    #10;

    a = 102;

    b = 154;

    cin = 0;

    #10;

    a = 82;

    b = 174;

    cin = 0;

    #10;

    a = 24;

    b = 231;

    cin = 1;

    #10;

    a = 199;

    b = 56;

    cin = 1;

    #10;

    a = 71;

    b = 184;

    cin = 1;

    #10;

    a = 64;

    b = 191;

    cin = 1;

    #10;

    a = 143;

    b = 113;

    cin = 0;

    #10;

    a = 239;

    b = 16;

    cin = 1;

    #10;

    a = 34;

    b = 221;

    cin = 1;

    #10;

    a = 157;

    b = 99;

    cin = 0;

    #10;

    a = 223;

    b = 33;

    cin = 0;

    #10;

    a = 172;

    b = 83;

    cin = 1;

    #10;

    a = 187;

    b = 69;

    cin = 0;

    #10;

    a = 150;

    b = 105;

    cin = 1;

    #10;

    a = 12;

    b = 244;

    cin = 0;

    #10;

    a = 241;

    b = 14;

    cin = 1;

    #10;

    a = 34;

    b = 222;

    cin = 0;

    #10;

    a = 180;

    b = 75;

    cin = 1;

    #10;

    a = 223;

    b = 33;

    cin = 0;

    #10;

    a = 122;

    b = 134;

    cin = 0;

    #10;

    a = 191;

    b = 65;

    cin = 0;

    #10;

    a = 252;

    b = 3;

    cin = 1;

    #10;

    a = 134;

    b = 122;

    cin = 0;

    #10;

    a = 71;

    b = 185;

    cin = 0;

    #10;

    a = 227;

    b = 28;

    cin = 1;

    #10;

    a = 70;

    b = 186;

    cin = 0;

    #10;

    a = 18;

    b = 237;

    cin = 1;

    #10;

    a = 154;

    b = 102;

    cin = 0;

    #10;

    a = 89;

    b = 167;

    cin = 0;

    #10;

    a = 154;

    b = 102;

    cin = 0;

    #10;

    a = 102;

    b = 154;

    cin = 0;

    #10;

    a = 205;

    b = 50;

    cin = 1;

    #10;

    a = 200;

    b = 56;

    cin = 0;

    #10;

    a = 186;

    b = 69;

    cin = 1;

    #10;

    a = 184;

    b = 71;

    cin = 1;

    #10;

    a = 186;

    b = 70;

    cin = 0;

    #10;

    a = 142;

    b = 113;

    cin = 1;

    #10;

    a = 39;

    b = 217;

    cin = 0;

    #10;

    a = 117;

    b = 138;

    cin = 1;

    #10;

    a = 127;

    b = 129;

    cin = 0;

    #10;

    a = 13;

    b = 242;

    cin = 1;

    #10;

    a = 224;

    b = 31;

    cin = 1;

    #10;

    a = 77;

    b = 178;

    cin = 1;

    #10;

    a = 142;

    b = 114;

    cin = 0;

    #10;

    a = 251;

    b = 5;

    cin = 0;

    #10;

    a = 114;

    b = 142;

    cin = 0;

    #10;

    a = 20;

    b = 235;

    cin = 1;

    #10;

    a = 209;

    b = 47;

    cin = 0;

    #10;

    a = 95;

    b = 161;

    cin = 0;

    #10;

    a = 32;

    b = 224;

    cin = 0;

    #10;

    a = 182;

    b = 74;

    cin = 0;

    #10;

    a = 98;

    b = 157;

    cin = 1;

    #10;

    a = 208;

    b = 48;

    cin = 0;

    #10;

    a = 107;

    b = 148;

    cin = 1;

    #10;

    a = 248;

    b = 8;

    cin = 0;

    #10;

    a = 190;

    b = 65;

    cin = 1;

    #10;

    a = 163;

    b = 93;

    cin = 0;

    #10;

    a = 23;

    b = 233;

    cin = 0;

    #10;

    a = 174;

    b = 82;

    cin = 0;

    #10;

    a = 86;

    b = 170;

    cin = 0;

    #10;

    a = 120;

    b = 135;

    cin = 1;

    #10;

    a = 187;

    b = 69;

    cin = 0;

    #10;

    a = 187;

    b = 68;

    cin = 1;

    #10;

    a = 135;

    b = 121;

    cin = 0;

    #10;

    a = 200;

    b = 56;

    cin = 0;

    #10;

    a = 126;

    b = 129;

    cin = 1;

    #10;

    a = 240;

    b = 16;

    cin = 0;

    #10;

    a = 216;

    b = 40;

    cin = 0;

    #10;

    a = 229;

    b = 27;

    cin = 0;

    #10;

    a = 239;

    b = 17;

    cin = 0;

    #10;

    a = 211;

    b = 45;

    cin = 0;

    #10;

    a = 157;

    b = 99;

    cin = 0;

    #10;

    a = 244;

    b = 12;

    cin = 0;

    #10;

    a = 253;

    b = 2;

    cin = 1;

    #10;

    a = 122;

    b = 134;

    cin = 0;

    #10;

    a = 12;

    b = 244;

    cin = 0;

    #10;

    a = 196;

    b = 59;

    cin = 1;

    #10;

    a = 39;

    b = 217;

    cin = 0;

    #10;

    a = 184;

    b = 72;

    cin = 0;

    #10;

    a = 207;

    b = 48;

    cin = 1;

    #10;

    a = 117;

    b = 139;

    cin = 0;

    #10;

    a = 85;

    b = 171;

    cin = 0;

    #10;

    a = 46;

    b = 209;

    cin = 1;

    #10;

    a = 40;

    b = 215;

    cin = 1;

    #10;

    a = 76;

    b = 179;

    cin = 1;

    #10;

    a = 17;

    b = 238;

    cin = 1;

    #10;

    a = 250;

    b = 6;

    cin = 0;

    #10;

    a = 201;

    b = 55;

    cin = 0;

    #10;

    a = 50;

    b = 205;

    cin = 1;

    #10;

    a = 35;

    b = 221;

    cin = 0;

    #10;

    a = 129;

    b = 126;

    cin = 1;

    #10;

    a = 72;

    b = 183;

    cin = 1;

    #10;

    a = 213;

    b = 43;

    cin = 0;

    #10;

    a = 20;

    b = 236;

    cin = 0;

    #10;

    a = 170;

    b = 86;

    cin = 0;

    #10;

    a = 171;

    b = 84;

    cin = 1;

    #10;

    a = 113;

    b = 142;

    cin = 1;

    #10;

    a = 243;

    b = 12;

    cin = 1;

    #10;

    a = 97;

    b = 159;

    cin = 0;

    #10;

    a = 149;

    b = 106;

    cin = 1;

    #10;

    a = 112;

    b = 143;

    cin = 1;

    #10;

    a = 114;

    b = 141;

    cin = 1;

    #10;

    a = 92;

    b = 163;

    cin = 1;

    #10;

    a = 81;

    b = 175;

    cin = 0;

    #10;

    a = 71;

    b = 184;

    cin = 1;

    #10;

    a = 187;

    b = 69;

    cin = 0;

    #10;

    a = 68;

    b = 187;

    cin = 1;

    #10;

    a = 147;

    b = 108;

    cin = 1;

    #10;

    a = 216;

    b = 39;

    cin = 1;

    #10;

    a = 235;

    b = 21;

    cin = 0;

    #10;

    a = 94;

    b = 161;

    cin = 1;

    #10;

    a = 34;

    b = 221;

    cin = 1;

    #10;

    a = 244;

    b = 12;

    cin = 0;

    #10;

    a = 253;

    b = 2;

    cin = 1;

    #10;

    a = 73;

    b = 183;

    cin = 0;

    #10;

    a = 91;

    b = 164;

    cin = 1;

    #10;

    a = 127;

    b = 129;

    cin = 0;

    #10;

    a = 122;

    b = 134;

    cin = 0;

    #10;

    a = 197;

    b = 58;

    cin = 1;

    #10;

    a = 9;

    b = 247;

    cin = 0;

    #10;

    a = 41;

    b = 215;

    cin = 0;

    #10;

    a = 216;

    b = 39;

    cin = 1;

    #10;

    a = 86;

    b = 169;

    cin = 1;

    #10;

    a = 42;

    b = 214;

    cin = 0;

    #10;

    a = 17;

    b = 238;

    cin = 1;

    #10;

    a = 246;

    b = 10;

    cin = 0;

    #10;

    a = 45;

    b = 211;

    cin = 0;

    #10;

    a = 252;

    b = 4;

    cin = 0;

    #10;

    a = 168;

    b = 88;

    cin = 0;

    #10;

    a = 231;

    b = 25;

    cin = 0;

    #10;

    a = 146;

    b = 110;

    cin = 0;

    #10;

    a = 156;

    b = 100;

    cin = 0;

    #10;

    a = 252;

    b = 4;

    cin = 0;

    #10;

    a = 85;

    b = 171;

    cin = 0;

    #10;

    a = 138;

    b = 118;

    cin = 0;

    #10;

    a = 79;

    b = 177;

    cin = 0;

    #10;

    a = 165;

    b = 90;

    cin = 1;

    #10;

    a = 160;

    b = 95;

    cin = 1;

    #10;

    a = 132;

    b = 124;

    cin = 0;

    #10;

    a = 56;

    b = 199;

    cin = 1;

    #10;

    a = 161;

    b = 95;

    cin = 0;

    #10;

    a = 1;

    b = 254;

    cin = 1;

    #10;

    a = 218;

    b = 37;

    cin = 1;

    #10;

    a = 91;

    b = 164;

    cin = 1;

    #10;

    a = 153;

    b = 103;

    cin = 0;

    #10;

    a = 158;

    b = 98;

    cin = 0;

    #10;

    a = 77;

    b = 179;

    cin = 0;

    #10;

    a = 115;

    b = 141;

    cin = 0;

    #10;

    a = 52;

    b = 204;

    cin = 0;

    #10;

    a = 82;

    b = 173;

    cin = 1;

    #10;

    a = 86;

    b = 170;

    cin = 0;

    #10;

    a = 32;

    b = 224;

    cin = 0;

    #10;

    a = 14;

    b = 242;

    cin = 0;

    #10;

    a = 87;

    b = 168;

    cin = 1;

    #10;

    a = 193;

    b = 62;

    cin = 1;

    #10;

    a = 218;

    b = 37;

    cin = 1;

    #10;

    a = 70;

    b = 186;

    cin = 0;

    #10;

    a = 206;

    b = 50;

    cin = 0;

    #10;

    a = 69;

    b = 186;

    cin = 1;

    #10;

    a = 52;

    b = 203;

    cin = 1;

    #10;

    a = 5;

    b = 250;

    cin = 1;

    #10;

    a = 116;

    b = 140;

    cin = 0;

    #10;

    a = 160;

    b = 95;

    cin = 1;

    #10;

    a = 196;

    b = 59;

    cin = 1;

    #10;

    a = 25;

    b = 231;

    cin = 0;

    #10;

    a = 141;

    b = 114;

    cin = 1;

    #10;

    a = 211;

    b = 44;

    cin = 1;

    #10;

    a = 203;

    b = 53;

    cin = 0;

    #10;

    a = 99;

    b = 156;

    cin = 1;

    #10;

    a = 154;

    b = 102;

    cin = 0;

    #10;

    a = 106;

    b = 149;

    cin = 1;

    #10;

    a = 133;

    b = 123;

    cin = 0;

    #10;

    a = 84;

    b = 171;

    cin = 1;

    #10;

    a = 142;

    b = 114;

    cin = 0;

    #10;

    a = 59;

    b = 197;

    cin = 0;

    #10;

    a = 17;

    b = 238;

    cin = 1;

    #10;

    a = 216;

    b = 39;

    cin = 1;

    #10;

    a = 202;

    b = 54;

    cin = 0;

    #10;

    a = 28;

    b = 227;

    cin = 1;

    #10;

    a = 83;

    b = 172;

    cin = 1;

    #10;

    a = 225;

    b = 30;

    cin = 1;

    #10;

    a = 192;

    b = 63;

    cin = 1;

    #10;

    a = 26;

    b = 229;

    cin = 1;

    #10;

    a = 240;

    b = 15;

    cin = 1;

    #10;

    a = 198;

    b = 58;

    cin = 0;

    #10;

    a = 206;

    b = 49;

    cin = 1;

    #10;

    a = 166;

    b = 90;

    cin = 0;

    #10;

    a = 180;

    b = 75;

    cin = 1;

    #10;

    a = 131;

    b = 125;

    cin = 0;

    #10;

    a = 218;

    b = 37;

    cin = 1;

    #10;

    a = 197;

    b = 59;

    cin = 0;

    #10;

    a = 138;

    b = 117;

    cin = 1;

    #10;

    a = 11;

    b = 245;

    cin = 0;

    #10;

    a = 7;

    b = 248;

    cin = 1;

    #10;

    a = 198;

    b = 58;

    cin = 0;

    #10;

    a = 135;

    b = 121;

    cin = 0;

    #10;

    a = 127;

    b = 128;

    cin = 1;

    #10;

    a = 85;

    b = 171;

    cin = 0;

    #10;

    a = 131;

    b = 124;

    cin = 1;

    #10;

    a = 219;

    b = 37;

    cin = 0;

    #10;

    a = 223;

    b = 33;

    cin = 0;

    #10;

    a = 164;

    b = 91;

    cin = 1;

    #10;

    a = 226;

    b = 29;

    cin = 1;

    #10;

    a = 160;

    b = 96;

    cin = 0;

    #10;

    a = 241;

    b = 15;

    cin = 0;

    #10;

    a = 48;

    b = 208;

    cin = 0;

    #10;

    a = 185;

    b = 70;

    cin = 1;

    #10;

    a = 110;

    b = 146;

    cin = 0;

    #10;

    a = 25;

    b = 231;

    cin = 0;

    #10;

    a = 80;

    b = 175;

    cin = 1;

    #10;

    a = 120;

    b = 136;

    cin = 0;

    #10;

    a = 141;

    b = 114;

    cin = 1;

    #10;

    a = 234;

    b = 21;

    cin = 1;

    #10;

    a = 44;

    b = 212;

    cin = 0;

    #10;

    a = 97;

    b = 158;

    cin = 1;

    #10;

    a = 92;

    b = 163;

    cin = 1;

    #10;

    a = 107;

    b = 148;

    cin = 1;

    #10;

    a = 78;

    b = 177;

    cin = 1;

    #10;

    a = 98;

    b = 158;

    cin = 0;

    #10;

    a = 77;

    b = 178;

    cin = 1;

    #10;

    a = 253;

    b = 3;

    cin = 0;

    #10;

    a = 210;

    b = 46;

    cin = 0;

    #10;

    a = 100;

    b = 156;

    cin = 0;

    #10;

    a = 44;

    b = 212;

    cin = 0;

    #10;

    a = 217;

    b = 39;

    cin = 0;

    #10;

    a = 48;

    b = 207;

    cin = 1;

    #10;

    a = 73;

    b = 183;

    cin = 0;

    #10;

    a = 88;

    b = 168;

    cin = 0;

    #10;

    a = 189;

    b = 67;

    cin = 0;

    #10;

    a = 112;

    b = 143;

    cin = 1;

    #10;

    a = 240;

    b = 15;

    cin = 1;

    #10;

    a = 32;

    b = 224;

    cin = 0;

    #10;

    a = 191;

    b = 65;

    cin = 0;

    #10;

    a = 61;

    b = 195;

    cin = 0;

    #10;

    a = 83;

    b = 172;

    cin = 1;

    #10;

    a = 18;

    b = 238;

    cin = 0;

    #10;

    a = 184;

    b = 71;

    cin = 1;

    #10;

    a = 143;

    b = 112;

    cin = 1;

    #10;

    a = 4;

    b = 252;

    cin = 0;

    #10;

    a = 150;

    b = 105;

    cin = 1;

    #10;

    a = 136;

    b = 120;

    cin = 0;

    #10;

    a = 191;

    b = 65;

    cin = 0;

    #10;

    a = 135;

    b = 120;

    cin = 1;

    #10;

    a = 78;

    b = 178;

    cin = 0;

    #10;

    a = 192;

    b = 64;

    cin = 0;

    #10;

    a = 147;

    b = 109;

    cin = 0;

    #10;

    a = 133;

    b = 122;

    cin = 1;

    #10;

    a = 64;

    b = 192;

    cin = 0;

    #10;

    a = 245;

    b = 10;

    cin = 1;

    #10;

    a = 200;

    b = 56;

    cin = 0;

    #10;

    a = 150;

    b = 106;

    cin = 0;

    #10;

    a = 12;

    b = 243;

    cin = 1;

    #10;

    a = 183;

    b = 73;

    cin = 0;

    #10;

    a = 173;

    b = 83;

    cin = 0;

    #10;

    a = 87;

    b = 169;

    cin = 0;

    #10;

    a = 122;

    b = 133;

    cin = 1;

    #10;

    a = 67;

    b = 189;

    cin = 0;

    #10;

    a = 254;

    b = 1;

    cin = 1;

    #10;

    a = 27;

    b = 229;

    cin = 0;

    #10;

    a = 232;

    b = 24;

    cin = 0;

    #10;

    a = 209;

    b = 46;

    cin = 1;

    #10;

    a = 145;

    b = 110;

    cin = 1;

    #10;

    a = 244;

    b = 11;

    cin = 1;

    #10;

    a = 158;

    b = 98;

    cin = 0;

    #10;

    a = 78;

    b = 178;

    cin = 0;

    #10;

    a = 161;

    b = 94;

    cin = 1;

    #10;

    a = 215;

    b = 41;

    cin = 0;

    #10;

    a = 163;

    b = 92;

    cin = 1;

    #10;

    a = 186;

    b = 70;

    cin = 0;

    #10;

    a = 225;

    b = 30;

    cin = 1;

    #10;

    a = 118;

    b = 137;

    cin = 1;

    #10;

    a = 57;

    b = 198;

    cin = 1;

    #10;

    a = 246;

    b = 10;

    cin = 0;

    #10;

    a = 21;

    b = 235;

    cin = 0;

    #10;

    a = 77;

    b = 179;

    cin = 0;

    #10;

    a = 18;

    b = 237;

    cin = 1;

    #10;

    a = 168;

    b = 87;

    cin = 1;

    #10;

    a = 177;

    b = 78;

    cin = 1;

    #10;

    a = 97;

    b = 159;

    cin = 0;

    #10;

    a = 127;

    b = 128;

    cin = 1;

    #10;

    a = 86;

    b = 169;

    cin = 1;

    #10;

    a = 182;

    b = 73;

    cin = 1;

    #10;

    a = 146;

    b = 109;

    cin = 1;

    #10;

    a = 251;

    b = 5;

    cin = 0;

    #10;

    a = 151;

    b = 105;

    cin = 0;

    #10;

    a = 8;

    b = 248;

    cin = 0;

    #10;

    a = 150;

    b = 105;

    cin = 1;

    #10;

    a = 119;

    b = 137;

    cin = 0;

    #10;

    a = 5;

    b = 250;

    cin = 1;

    #10;

    a = 140;

    b = 116;

    cin = 0;

    #10;

    a = 8;

    b = 248;

    cin = 0;

    #10;

    a = 211;

    b = 44;

    cin = 1;

    #10;

    a = 26;

    b = 230;

    cin = 0;

    #10;

    a = 42;

    b = 214;

    cin = 0;

    #10;

    a = 230;

    b = 26;

    cin = 0;

    #10;

    a = 240;

    b = 15;

    cin = 1;

    #10;

    a = 73;

    b = 183;

    cin = 0;

    #10;

    a = 240;

    b = 16;

    cin = 0;

    #10;

    a = 212;

    b = 44;

    cin = 0;

    #10;

    a = 163;

    b = 92;

    cin = 1;

    #10;

    a = 168;

    b = 88;

    cin = 0;

    #10;

    a = 150;

    b = 105;

    cin = 1;

    #10;

    a = 239;

    b = 17;

    cin = 0;

    #10;

    a = 37;

    b = 219;

    cin = 0;

    #10;

    a = 191;

    b = 64;

    cin = 1;

    #10;

    a = 227;

    b = 28;

    cin = 1;

    #10;

    a = 137;

    b = 118;

    cin = 1;

    #10;

    a = 132;

    b = 123;

    cin = 1;

    #10;

    a = 244;

    b = 12;

    cin = 0;

    #10;

    a = 102;

    b = 153;

    cin = 1;

    #10;

    a = 204;

    b = 52;

    cin = 0;

    #10;

    a = 6;

    b = 250;

    cin = 0;

    #10;

    a = 240;

    b = 15;

    cin = 1;

    #10;

    a = 126;

    b = 129;

    cin = 1;

    #10;

    a = 131;

    b = 124;

    cin = 1;

    #10;

    a = 49;

    b = 207;

    cin = 0;

    #10;

    a = 234;

    b = 22;

    cin = 0;

    #10;

    a = 38;

    b = 217;

    cin = 1;

    #10;

    a = 102;

    b = 153;

    cin = 1;

    #10;

    a = 161;

    b = 95;

    cin = 0;

    #10;

    a = 218;

    b = 38;

    cin = 0;

    #10;

    a = 95;

    b = 160;

    cin = 1;

    #10;

    a = 79;

    b = 176;

    cin = 1;

    #10;

    a = 50;

    b = 206;

    cin = 0;

    #10;

    a = 141;

    b = 115;

    cin = 0;

    #10;

    a = 14;

    b = 242;

    cin = 0;

    #10;

    a = 36;

    b = 219;

    cin = 1;

    #10;

    a = 89;

    b = 167;

    cin = 0;

    #10;

    a = 70;

    b = 185;

    cin = 1;

    #10;

    a = 253;

    b = 2;

    cin = 1;

    #10;

    a = 170;

    b = 86;

    cin = 0;

    #10;

    a = 178;

    b = 77;

    cin = 1;

    #10;

    a = 192;

    b = 64;

    cin = 0;

    #10;

    a = 204;

    b = 51;

    cin = 1;

    #10;

    a = 57;

    b = 199;

    cin = 0;

    #10;

    a = 246;

    b = 10;

    cin = 0;

    #10;

    a = 110;

    b = 145;

    cin = 1;

    #10;

    a = 123;

    b = 133;

    cin = 0;

    #10;

    a = 182;

    b = 74;

    cin = 0;

    #10;

    a = 106;

    b = 149;

    cin = 1;

    #10;

    a = 229;

    b = 27;

    cin = 0;

    #10;

    a = 238;

    b = 18;

    cin = 0;

    #10;

    a = 156;

    b = 100;

    cin = 0;

    #10;

    a = 56;

    b = 199;

    cin = 1;

    #10;

    a = 193;

    b = 62;

    cin = 1;

    #10;

    a = 140;

    b = 115;

    cin = 1;

    #10;

    a = 210;

    b = 46;

    cin = 0;

    #10;

    a = 252;

    b = 4;

    cin = 0;

    #10;

    a = 51;

    b = 204;

    cin = 1;

    #10;

    a = 253;

    b = 3;

    cin = 0;

    #10;

    a = 201;

    b = 55;

    cin = 0;

    #10;

    a = 152;

    b = 103;

    cin = 1;

    #10;

    a = 142;

    b = 113;

    cin = 1;

    #10;

    a = 231;

    b = 25;

    cin = 0;

    #10;

    a = 10;

    b = 246;

    cin = 0;

    #10;

    a = 194;

    b = 61;

    cin = 1;

    #10;

    a = 222;

    b = 34;

    cin = 0;

    #10;

    a = 11;

    b = 245;

    cin = 0;

    #10;

    a = 147;

    b = 108;

    cin = 1;

    #10;

    a = 208;

    b = 48;

    cin = 0;

    #10;

    a = 49;

    b = 206;

    cin = 1;

    #10;

    a = 0;

    b = 255;

    cin = 1;

    #10;

    a = 92;

    b = 163;

    cin = 1;

    #10;

    a = 213;

    b = 42;

    cin = 1;

    #10;

    a = 56;

    b = 200;

    cin = 0;

    #10;

    a = 84;

    b = 171;

    cin = 1;

    #10;

    a = 172;

    b = 83;

    cin = 1;

    #10;

    a = 245;

    b = 10;

    cin = 1;

    #10;

    a = 96;

    b = 159;

    cin = 1;

    #10;

    a = 208;

    b = 48;

    cin = 0;

    #10;

    a = 148;

    b = 108;

    cin = 0;

    #10;

    a = 142;

    b = 114;

    cin = 0;

    #10;

    a = 39;

    b = 217;

    cin = 0;

    #10;

    a = 231;

    b = 25;

    cin = 0;

    #10;

    a = 206;

    b = 49;

    cin = 1;

    #10;

    a = 237;

    b = 18;

    cin = 1;

    #10;

    a = 183;

    b = 73;

    cin = 0;

    #10;

    a = 124;

    b = 131;

    cin = 1;

    #10;

    a = 167;

    b = 89;

    cin = 0;

    #10;

    a = 151;

    b = 105;

    cin = 0;

    #10;

    a = 19;

    b = 237;

    cin = 0;

    #10;

    a = 212;

    b = 44;

    cin = 0;

    #10;

    a = 234;

    b = 22;

    cin = 0;

    #10;

    a = 19;

    b = 236;

    cin = 1;

    #10;

    a = 169;

    b = 87;

    cin = 0;

    #10;

    a = 106;

    b = 150;

    cin = 0;

    #10;

    a = 251;

    b = 5;

    cin = 0;

    #10;

    a = 108;

    b = 148;

    cin = 0;

    #10;

    a = 190;

    b = 65;

    cin = 1;

    #10;

    a = 81;

    b = 174;

    cin = 1;

    #10;

    a = 134;

    b = 121;

    cin = 1;

    #10;

    a = 209;

    b = 47;

    cin = 0;

    #10;

    a = 203;

    b = 53;

    cin = 0;

    #10;

    a = 8;

    b = 248;

    cin = 0;

    #10;

    a = 247;

    b = 8;

    cin = 1;

    #10;

    a = 189;

    b = 67;

    cin = 0;

    #10;

    a = 72;

    b = 184;

    cin = 0;

    #10;

    a = 179;

    b = 76;

    cin = 1;

    #10;

    a = 250;

    b = 5;

    cin = 1;

    #10;

    a = 231;

    b = 25;

    cin = 0;

    #10;

    a = 54;

    b = 201;

    cin = 1;

    #10;

    a = 43;

    b = 212;

    cin = 1;

    #10;

    a = 83;

    b = 173;

    cin = 0;

    #10;

    a = 33;

    b = 223;

    cin = 0;

    #10;

    a = 31;

    b = 225;

    cin = 0;

    #10;

    a = 45;

    b = 211;

    cin = 0;

    #10;

    a = 7;

    b = 248;

    cin = 1;

    #10;

    a = 165;

    b = 90;

    cin = 1;

    #10;

    a = 61;

    b = 194;

    cin = 1;

    #10;

    a = 158;

    b = 97;

    cin = 1;

    #10;

    a = 158;

    b = 97;

    cin = 1;

    #10;

    a = 184;

    b = 72;

    cin = 0;

    #10;

    a = 62;

    b = 194;

    cin = 0;

    #10;

    a = 255;

    b = 1;

    cin = 0;

    #10;

    a = 160;

    b = 96;

    cin = 0;

    #10;

    a = 117;

    b = 139;

    cin = 0;

    #10;

    a = 210;

    b = 45;

    cin = 1;

    #10;

    a = 44;

    b = 211;

    cin = 1;

    #10;

    a = 117;

    b = 139;

    cin = 0;

    #10;

    a = 90;

    b = 166;

    cin = 0;

    #10;

    a = 51;

    b = 204;

    cin = 1;

    #10;

    a = 75;

    b = 180;

    cin = 1;

    #10;

    a = 234;

    b = 21;

    cin = 1;

    #10;

    a = 188;

    b = 67;

    cin = 1;

    #10;

    a = 105;

    b = 151;

    cin = 0;

    #10;

    a = 16;

    b = 239;

    cin = 1;

    #10;

    a = 126;

    b = 130;

    cin = 0;

    #10;

    a = 141;

    b = 114;

    cin = 1;

    #10;

    a = 201;

    b = 55;

    cin = 0;

    #10;

    a = 183;

    b = 72;

    cin = 1;

    #10;

    a = 71;

    b = 184;

    cin = 1;

    #10;

    a = 49;

    b = 207;

    cin = 0;

    #10;

    a = 76;

    b = 180;

    cin = 0;

    #10;

    a = 65;

    b = 191;

    cin = 0;

    #10;

    a = 82;

    b = 173;

    cin = 1;

    #10;

    a = 110;

    b = 145;

    cin = 1;

    #10;

    a = 54;

    b = 201;

    cin = 1;

    #10;

    a = 161;

    b = 94;

    cin = 1;

    #10;

    a = 13;

    b = 243;

    cin = 0;

    #10;

    a = 236;

    b = 20;

    cin = 0;

    #10;

    a = 217;

    b = 39;

    cin = 0;

    #10;

    a = 217;

    b = 39;

    cin = 0;

    #10;

    a = 70;

    b = 185;

    cin = 1;

    #10;

    a = 36;

    b = 220;

    cin = 0;

    #10;

    a = 171;

    b = 84;

    cin = 1;

    #10;

    a = 83;

    b = 172;

    cin = 1;

    #10;

    a = 6;

    b = 250;

    cin = 0;

    #10;

    a = 182;

    b = 74;

    cin = 0;

    #10;

    a = 62;

    b = 193;

    cin = 1;

    #10;

    a = 211;

    b = 44;

    cin = 1;

    #10;

    a = 79;

    b = 177;

    cin = 0;

    #10;

    a = 164;

    b = 91;

    cin = 1;

    #10;

    a = 168;

    b = 88;

    cin = 0;

    #10;

    a = 123;

    b = 133;

    cin = 0;

    #10;

    a = 147;

    b = 109;

    cin = 0;

    #10;

    a = 4;

    b = 252;

    cin = 0;

    #10;

    a = 45;

    b = 210;

    cin = 1;

    #10;

    a = 1;

    b = 255;

    cin = 0;

    #10;

    a = 85;

    b = 171;

    cin = 0;

    #10;

    a = 53;

    b = 202;

    cin = 1;

    #10;

    a = 68;

    b = 188;

    cin = 0;

    #10;

    a = 144;

    b = 112;

    cin = 0;

    #10;

    a = 131;

    b = 125;

    cin = 0;

    #10;

    a = 190;

    b = 66;

    cin = 0;

    #10;

    a = 149;

    b = 107;

    cin = 0;

    #10;

    a = 236;

    b = 20;

    cin = 0;

    #10;

    a = 235;

    b = 20;

    cin = 1;

    #10;

    a = 7;

    b = 248;

    cin = 1;

    #10;

    a = 57;

    b = 199;

    cin = 0;

    #10;

    a = 2;

    b = 254;

    cin = 0;

    #10;

    a = 163;

    b = 93;

    cin = 0;

    #10;

    a = 223;

    b = 32;

    cin = 1;

    #10;

    a = 1;

    b = 255;

    cin = 0;

    #10;

    a = 121;

    b = 134;

    cin = 1;

    #10;

    a = 58;

    b = 198;

    cin = 0;

    #10;

    a = 59;

    b = 197;

    cin = 0;

    #10;

    a = 238;

    b = 18;

    cin = 0;

    #10;

    a = 21;

    b = 235;

    cin = 0;

    #10;

    a = 74;

    b = 181;

    cin = 1;

    #10;

    a = 130;

    b = 126;

    cin = 0;

    #10;

    a = 197;

    b = 59;

    cin = 0;

    #10;

    a = 118;

    b = 138;

    cin = 0;

    #10;

    a = 103;

    b = 153;

    cin = 0;

    #10;

    a = 105;

    b = 151;

    cin = 0;

    #10;

    a = 236;

    b = 19;

    cin = 1;

    #10;

    a = 39;

    b = 216;

    cin = 1;

    #10;

    a = 12;

    b = 244;

    cin = 0;

    #10;

    a = 8;

    b = 248;

    cin = 0;

    #10;

    a = 125;

    b = 131;

    cin = 0;

    #10;

    a = 242;

    b = 13;

    cin = 1;

    #10;

    a = 240;

    b = 15;

    cin = 1;

    #10;

    a = 121;

    b = 135;

    cin = 0;

    #10;

    a = 11;

    b = 244;

    cin = 1;

    #10;

    a = 150;

    b = 105;

    cin = 1;

    #10;

    a = 154;

    b = 101;

    cin = 1;

    #10;

    a = 226;

    b = 30;

    cin = 0;

    #10;

    a = 74;

    b = 181;

    cin = 1;

    #10;

    a = 240;

    b = 15;

    cin = 1;

    #10;

    a = 186;

    b = 69;

    cin = 1;

    #10;

    a = 117;

    b = 139;

    cin = 0;

    #10;

    a = 157;

    b = 98;

    cin = 1;

    #10;

    a = 224;

    b = 31;

    cin = 1;

    #10;

    a = 2;

    b = 254;

    cin = 0;

    #10;

    a = 84;

    b = 171;

    cin = 1;

    #10;

    a = 174;

    b = 81;

    cin = 1;

    #10;

    a = 121;

    b = 134;

    cin = 1;

    #10;

    a = 164;

    b = 91;

    cin = 1;

    #10;

    a = 228;

    b = 27;

    cin = 1;

    #10;

    a = 228;

    b = 27;

    cin = 1;

    #10;

    a = 145;

    b = 110;

    cin = 1;

    #10;

    a = 104;

    b = 152;

    cin = 0;

    #10;

    a = 113;

    b = 142;

    cin = 1;

    #10;

    a = 206;

    b = 49;

    cin = 1;

    #10;

    a = 174;

    b = 82;

    cin = 0;

    #10;

    a = 187;

    b = 68;

    cin = 1;

    #10;

    a = 182;

    b = 74;

    cin = 0;

    #10;

    a = 67;

    b = 188;

    cin = 1;

    #10;

    a = 146;

    b = 109;

    cin = 1;

    #10;

    a = 154;

    b = 102;

    cin = 0;

    #10;

    a = 48;

    b = 207;

    cin = 1;

    #10;

    a = 102;

    b = 154;

    cin = 0;

    #10;

    a = 26;

    b = 230;

    cin = 0;

    #10;

    a = 224;

    b = 31;

    cin = 1;

    #10;

    a = 121;

    b = 135;

    cin = 0;

    #10;

    a = 249;

    b = 6;

    cin = 1;

    #10;

    a = 21;

    b = 234;

    cin = 1;

    #10;

    a = 180;

    b = 76;

    cin = 0;

    #10;

    a = 115;

    b = 141;

    cin = 0;

    #10;

    a = 114;

    b = 142;

    cin = 0;

    #10;

    a = 118;

    b = 138;

    cin = 0;

    #10;

    a = 236;

    b = 20;

    cin = 0;

    #10;

    a = 53;

    b = 202;

    cin = 1;

    #10;

    a = 205;

    b = 51;

    cin = 0;

    #10;

    a = 88;

    b = 168;

    cin = 0;

    #10;

    a = 33;

    b = 222;

    cin = 1;

    #10;

    a = 7;

    b = 249;

    cin = 0;

    #10;

    a = 87;

    b = 169;

    cin = 0;

    #10;

    a = 205;

    b = 50;

    cin = 1;

    #10;

    a = 234;

    b = 21;

    cin = 1;

    #10;

    a = 240;

    b = 16;

    cin = 0;

    #10;

    a = 35;

    b = 221;

    cin = 0;

    #10;

    a = 255;

    b = 0;

    cin = 1;

    #10;

    a = 147;

    b = 109;

    cin = 0;

    #10;

    a = 236;

    b = 19;

    cin = 1;

    #10;

    a = 189;

    b = 67;

    cin = 0;

    #10;

    a = 172;

    b = 84;

    cin = 0;

    #10;

    a = 210;

    b = 45;

    cin = 1;

    #10;

    a = 190;

    b = 65;

    cin = 1;

    #10;

    a = 99;

    b = 157;

    cin = 0;

    #10;

    a = 171;

    b = 85;

    cin = 0;

    #10;

    a = 227;

    b = 28;

    cin = 1;

    #10;

    a = 141;

    b = 114;

    cin = 1;

    #10;

    a = 234;

    b = 22;

    cin = 0;

    #10;

    a = 34;

    b = 222;

    cin = 0;

    #10;

    a = 241;

    b = 15;

    cin = 0;

    #10;

    a = 80;

    b = 175;

    cin = 1;

    #10;

    a = 210;

    b = 46;

    cin = 0;

    #10;

    a = 47;

    b = 209;

    cin = 0;

    #10;

    a = 97;

    b = 159;

    cin = 0;

    #10;

    a = 136;

    b = 120;

    cin = 0;

    #10;

    a = 242;

    b = 13;

    cin = 1;

    #10;

    a = 239;

    b = 16;

    cin = 1;

    #10;

    a = 254;

    b = 2;

    cin = 0;

    #10;

    a = 107;

    b = 148;

    cin = 1;

    #10;

    a = 34;

    b = 221;

    cin = 1;

    #10;

    a = 16;

    b = 240;

    cin = 0;

    #10;

    a = 50;

    b = 205;

    cin = 1;

    #10;

    a = 141;

    b = 115;

    cin = 0;

    #10;

    a = 248;

    b = 8;

    cin = 0;

    #10;

    a = 121;

    b = 135;

    cin = 0;

    #10;

    a = 31;

    b = 225;

    cin = 0;

    #10;

    a = 199;

    b = 57;

    cin = 0;

    #10;

    a = 72;

    b = 184;

    cin = 0;

    #10;

    a = 13;

    b = 243;

    cin = 0;

    #10;

    a = 205;

    b = 51;

    cin = 0;

    #10;

    a = 69;

    b = 186;

    cin = 1;

    #10;

    a = 122;

    b = 133;

    cin = 1;

    #10;

    a = 57;

    b = 198;

    cin = 1;

    #10;

    a = 59;

    b = 197;

    cin = 0;

    #10;

    a = 78;

    b = 177;

    cin = 1;

    #10;

    a = 195;

    b = 61;

    cin = 0;

    #10;

    a = 78;

    b = 177;

    cin = 1;

    #10;

    a = 100;

    b = 156;

    cin = 0;

    #10;

    a = 100;

    b = 156;

    cin = 0;

    #10;

    a = 144;

    b = 111;

    cin = 1;

    #10;

    a = 82;

    b = 174;

    cin = 0;

    #10;

    a = 153;

    b = 102;

    cin = 1;

    #10;

    a = 55;

    b = 200;

    cin = 1;

    #10;

    a = 125;

    b = 131;

    cin = 0;

    #10;

    a = 181;

    b = 75;

    cin = 0;

    #10;

    a = 22;

    b = 234;

    cin = 0;

    #10;

    a = 246;

    b = 10;

    cin = 0;

    #10;

    a = 183;

    b = 73;

    cin = 0;

    #10;

    a = 238;

    b = 17;

    cin = 1;

    #10;

    a = 222;

    b = 33;

    cin = 1;

    #10;

    a = 112;

    b = 143;

    cin = 1;

    #10;

    a = 36;

    b = 219;

    cin = 1;

    #10;

    a = 4;

    b = 252;

    cin = 0;

    #10;

    a = 158;

    b = 98;

    cin = 0;

    #10;

    a = 91;

    b = 165;

    cin = 0;

    #10;

    a = 121;

    b = 134;

    cin = 1;

    #10;

    a = 166;

    b = 90;

    cin = 0;

    #10;

    a = 254;

    b = 1;

    cin = 1;

    #10;

    a = 173;

    b = 83;

    cin = 0;

    #10;

    a = 98;

    b = 158;

    cin = 0;

    #10;

    a = 39;

    b = 216;

    cin = 1;

    #10;

    a = 7;

    b = 249;

    cin = 0;

    #10;

    a = 77;

    b = 179;

    cin = 0;

    #10;

    a = 51;

    b = 204;

    cin = 1;

    #10;

    a = 118;

    b = 138;

    cin = 0;

    #10;

    a = 165;

    b = 91;

    cin = 0;

    #10;

    a = 58;

    b = 198;

    cin = 0;

    #10;

    a = 43;

    b = 212;

    cin = 1;

    #10;

    a = 142;

    b = 114;

    cin = 0;

    #10;

    a = 33;

    b = 223;

    cin = 0;

    #10;

    a = 231;

    b = 24;

    cin = 1;

    #10;

    a = 49;

    b = 206;

    cin = 1;

    #10;

    a = 44;

    b = 211;

    cin = 1;

    #10;

    a = 159;

    b = 96;

    cin = 1;

    #10;

    a = 12;

    b = 243;

    cin = 1;

    #10;

    a = 120;

    b = 135;

    cin = 1;

    #10;

    a = 162;

    b = 94;

    cin = 0;

    #10;

    a = 197;

    b = 59;

    cin = 0;

    #10;

    a = 208;

    b = 48;

    cin = 0;

    #10;

    a = 185;

    b = 70;

    cin = 1;

    #10;

    a = 99;

    b = 156;

    cin = 1;

    #10;

    a = 50;

    b = 205;

    cin = 1;

    #10;

    a = 103;

    b = 152;

    cin = 1;

    #10;

    a = 73;

    b = 182;

    cin = 1;

    #10;

    a = 101;

    b = 155;

    cin = 0;

    #10;

    a = 72;

    b = 184;

    cin = 0;

    #10;

    a = 238;

    b = 17;

    cin = 1;

    #10;

    a = 169;

    b = 86;

    cin = 1;

    #10;

    a = 238;

    b = 18;

    cin = 0;

    #10;

    a = 244;

    b = 12;

    cin = 0;

    #10;

    a = 137;

    b = 119;

    cin = 0;

    #10;

    a = 130;

    b = 125;

    cin = 1;

    #10;

    a = 250;

    b = 5;

    cin = 1;

    #10;

    a = 202;

    b = 53;

    cin = 1;

    #10;

    a = 78;

    b = 178;

    cin = 0;

    #10;

    a = 199;

    b = 57;

    cin = 0;

    #10;

    a = 235;

    b = 20;

    cin = 1;

    #10;

    a = 117;

    b = 138;

    cin = 1;

    #10;

    a = 45;

    b = 211;

    cin = 0;

    #10;

    a = 14;

    b = 241;

    cin = 1;

    #10;

    a = 175;

    b = 80;

    cin = 1;

    #10;

    a = 153;

    b = 102;

    cin = 1;

    #10;

    a = 119;

    b = 137;

    cin = 0;

    #10;

    a = 30;

    b = 226;

    cin = 0;

    #10;

    a = 125;

    b = 131;

    cin = 0;

    #10;

    a = 85;

    b = 171;

    cin = 0;

    #10;

    a = 206;

    b = 50;

    cin = 0;

    #10;

    a = 94;

    b = 162;

    cin = 0;

    #10;

    a = 234;

    b = 22;

    cin = 0;

    #10;

    a = 212;

    b = 43;

    cin = 1;

    #10;

    a = 122;

    b = 133;

    cin = 1;

    #10;

    a = 77;

    b = 178;

    cin = 1;

    #10;

    a = 96;

    b = 159;

    cin = 1;

    #10;

    a = 212;

    b = 43;

    cin = 1;

    #10;

    a = 181;

    b = 74;

    cin = 1;

    #10;

    a = 164;

    b = 91;

    cin = 1;

    #10;

    a = 233;

    b = 23;

    cin = 0;

    #10;

    a = 115;

    b = 141;

    cin = 0;

    #10;

    a = 237;

    b = 18;

    cin = 1;

    #10;

    a = 149;

    b = 106;

    cin = 1;

    #10;

    a = 150;

    b = 106;

    cin = 0;

    #10;

    a = 202;

    b = 53;

    cin = 1;

    #10;

    a = 168;

    b = 87;

    cin = 1;

    #10;

    a = 25;

    b = 231;

    cin = 0;

    #10;

    a = 173;

    b = 83;

    cin = 0;

    #10;

    a = 232;

    b = 24;

    cin = 0;

    #10;

    a = 131;

    b = 124;

    cin = 1;

    #10;

    a = 180;

    b = 75;

    cin = 1;

    #10;

    a = 70;

    b = 186;

    cin = 0;

    #10;

    a = 22;

    b = 233;

    cin = 1;

    #10;

    a = 233;

    b = 23;

    cin = 0;

    #10;

    a = 202;

    b = 54;

    cin = 0;

    #10;

    a = 12;

    b = 243;

    cin = 1;

    #10;

    a = 99;

    b = 157;

    cin = 0;

    #10;

    a = 87;

    b = 169;

    cin = 0;

    #10;

    a = 3;

    b = 253;

    cin = 0;

    #10;

    a = 190;

    b = 65;

    cin = 1;

    #10;

    a = 175;

    b = 80;

    cin = 1;

    #10;

    a = 197;

    b = 58;

    cin = 1;

    #10;

    a = 212;

    b = 43;

    cin = 1;

    #10;

    a = 151;

    b = 104;

    cin = 1;

    #10;

    a = 76;

    b = 180;

    cin = 0;

    #10;

    a = 50;

    b = 206;

    cin = 0;

    #10;

    a = 187;

    b = 69;

    cin = 0;

    #10;

    a = 147;

    b = 109;

    cin = 0;

    #10;

    a = 238;

    b = 17;

    cin = 1;

    #10;

    a = 191;

    b = 65;

    cin = 0;

    #10;

    a = 82;

    b = 173;

    cin = 1;

    #10;

    a = 205;

    b = 51;

    cin = 0;

    #10;

    a = 216;

    b = 39;

    cin = 1;

    #10;

    a = 27;

    b = 228;

    cin = 1;

    #10;

    a = 189;

    b = 66;

    cin = 1;

    #10;

    a = 234;

    b = 22;

    cin = 0;

    #10;

    a = 51;

    b = 205;

    cin = 0;

    #10;

    a = 21;

    b = 235;

    cin = 0;

    #10;

    a = 52;

    b = 204;

    cin = 0;

    #10;

    a = 174;

    b = 82;

    cin = 0;

    #10;

    a = 56;

    b = 200;

    cin = 0;

    #10;

    a = 27;

    b = 229;

    cin = 0;

    #10;

    a = 94;

    b = 162;

    cin = 0;

    #10;

    a = 80;

    b = 175;

    cin = 1;

    #10;

    a = 87;

    b = 168;

    cin = 1;

    #10;

    a = 87;

    b = 168;

    cin = 1;

    #10;

    a = 232;

    b = 23;

    cin = 1;

    #10;

    a = 152;

    b = 103;

    cin = 1;

    #10;

    a = 226;

    b = 30;

    cin = 0;

    #10;

    a = 208;

    b = 47;

    cin = 1;

    #10;

    a = 75;

    b = 181;

    cin = 0;

    #10;

    a = 159;

    b = 96;

    cin = 1;

    #10;

    a = 162;

    b = 93;

    cin = 1;

    #10;

    a = 125;

    b = 130;

    cin = 1;

    #10;

    a = 229;

    b = 27;

    cin = 0;

    #10;

    a = 133;

    b = 122;

    cin = 1;

    #10;

    a = 47;

    b = 208;

    cin = 1;

    #10;

    a = 187;

    b = 69;

    cin = 0;

    #10;

    a = 242;

    b = 14;

    cin = 0;

    #10;

    a = 86;

    b = 170;

    cin = 0;

    #10;

    a = 119;

    b = 136;

    cin = 1;

    #10;

    a = 253;

    b = 3;

    cin = 0;

    #10;

    a = 14;

    b = 241;

    cin = 1;

    #10;

    a = 90;

    b = 165;

    cin = 1;

    #10;

    a = 29;

    b = 226;

    cin = 1;

    #10;

    a = 168;

    b = 87;

    cin = 1;

    #10;

    a = 220;

    b = 36;

    cin = 0;

    #10;

    a = 74;

    b = 182;

    cin = 0;

    #10;

    a = 231;

    b = 25;

    cin = 0;

    #10;

    a = 86;

    b = 169;

    cin = 1;

    #10;

    a = 226;

    b = 30;

    cin = 0;

    #10;

    a = 19;

    b = 237;

    cin = 0;

    #10;

    a = 87;

    b = 169;

    cin = 0;

    #10;

    a = 226;

    b = 29;

    cin = 1;

    #10;

    a = 175;

    b = 80;

    cin = 1;

    #10;

    #50;

    $finish;
  end
endmodule
