//gets the packet from generator and drive the transaction paket items into interface (interface is connected to DUT, so the items driven into interface signal will get driven in to DUT) 

class driver;

    //used to count the number of transactions
    int no_transactions;

    //creating virtual interface handle
    virtual vendingmachine_intf vendingmachine_vif;

    //creating mailbox handle
    mailbox gen2driv;

    //constructor
    function new(virtual vendingmachine_intf vendingmachine_vif,mailbox gen2driv);
        //getting the interface
        this.vendingmachine_vif = vendingmachine_vif;
        //getting the mailbox handles from  environment 
        this.gen2driv = gen2driv;
    endfunction

    //Reset task, Reset the Interface signals to default/initial values
    task reset;
        wait(vendingmachine_vif.rst);
        $display("--------- [DRIVER] Reset Started ---------");
        wait(!vendingmachine_vif.rst);
        $display("--------- [DRIVER] Reset Ended ---------");
    endtask

    //drivers the transaction items to interface signals
    task drive;
        transaction trans;
        gen2driv.get(trans);
        vendingmachine_vif.coin_in=trans.coin_in;
        vendingmachine_vif.button_in=trans.button_in;
        no_transactions++;
        @(posedge vendingmachine_vif.clk);
    endtask


    task main;
        wait(!vendingmachine_vif.rst);
        forever
            drive();
   endtask

endclass
