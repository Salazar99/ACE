`timescale 1ns/1ns

module test;

  logic clk;

  logic [2:0] A;

  logic [2:0] B;

  logic A_greater;

  logic A_equal;

  logic A_less;


  // Device Under Test (DUT)

  comparator_3bit dut(
    .clk(clk),
    .A(A),
    .B(B),
    .A_greater(A_greater),
    .A_equal(A_equal),
    .A_less(A_less)
  );


  always #5 clk = ~clk;


  initial begin

    $dumpfile("comparator_3bit.vcd");

    $dumpvars(0, test);

    clk = 0;

    A = 0;

    B = 0;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 3;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 6;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 1;

    B = 0;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 5;

    B = 3;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 6;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 7;

    B = 2;

    #10;

    A = 0;

    B = 2;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 1;

    B = 3;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 1;

    B = 4;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 3;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 1;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 3;

    B = 1;

    #10;

    A = 3;

    B = 6;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 7;

    B = 1;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 6;

    B = 0;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 0;

    B = 1;

    #10;

    A = 2;

    B = 7;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 1;

    B = 2;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 5;

    B = 1;

    #10;

    A = 0;

    B = 4;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 1;

    B = 6;

    #10;

    A = 5;

    B = 7;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 4;

    B = 1;

    #10;

    A = 4;

    B = 0;

    #10;

    A = 5;

    B = 4;

    #10;

    A = 2;

    B = 0;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 0;

    B = 7;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 0;

    B = 3;

    #10;

    A = 7;

    B = 4;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 2;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 7;

    B = 3;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 2;

    B = 1;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 5;

    B = 2;

    #10;

    A = 2;

    B = 4;

    #10;

    A = 6;

    B = 4;

    #10;

    A = 2;

    B = 5;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 2;

    B = 6;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 4;

    B = 7;

    #10;

    A = 3;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 1;

    B = 5;

    #10;

    A = 3;

    B = 2;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 5;

    B = 0;

    #10;

    A = 6;

    B = 5;

    #10;

    A = 3;

    B = 0;

    #10;

    A = 0;

    B = 6;

    #10;

    A = 4;

    B = 3;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 5;

    B = 6;

    #10;

    A = 7;

    B = 5;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 1;

    #10;

    A = 6;

    B = 7;

    #10;

    A = 3;

    B = 7;

    #10;

    A = 3;

    B = 4;

    #10;

    A = 4;

    B = 2;

    #10;

    A = 7;

    B = 0;

    #10;

    A = 4;

    B = 5;

    #10;

    A = 0;

    B = 5;

    #10;

    A = 5;

    B = 4;

    #10;

    #50;

    $finish;
  end
endmodule
